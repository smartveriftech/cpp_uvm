// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
PH+KUF.HEK.GL0*TZ*#NJ1,M4(5/6L DF\;3Z:WQPING?</<**P'_O-)UABUT%/+,
P 3T\+_[/A/D6X+E[V>XW9L$?>!1R*=QHFIB-4>/Y""\<G7EK->=G-;[9P=:QHT#I
P3>7*M\+QN\JNPZ*W\_A(_5Z8FHBSZH*^=5A^Z;Q;\X1@O7-;9<D<J1(NUSB(T=[W
P*NR$P$38K*"/.*R""Q@3JH?_L!V+#<TE/(XBMZ>UXGD1A63@OJD6>FT".%(4H;[1
P+8A^^3Z'2!-/WQ-:RCY/-W?T$+$G4_$5UHYBZHJMHPT]W<72-M8@6 ]6UGI4WN)2
`endprotected128

