// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Guard to prevent multiple inclusions
`protected128
P)D=136R:<P_MF(WW 2;=7#3I7B5L#A.>I?PH&V\R1(<_UU.-)M!A&W&]WM03N5,&
PT73Q(X74\]_:X9%5X@L;R/J?Z,M?[F+&-J/ BC[N>!_61D*G=^Z'K<,B7A178L%?
PW;24P@^E4,4\!07'G2.=[AA6]&.6Z**I%[$41+0-@>6-CPSZRCOD( =;XL]$;-K:
P3O>>N1H?<%-=[X!#96@)<<KX((Y5:HUT($[$8^0OJJEM(=:1B0K@X67("_TD*E\4
PF(\BQI5Y5R@A>EL)/@:A8V)9B$TGV@UV,;E8KM!B3Z)1:91GK@ -:,C#D="YV7W,
P:>2A:HXE=&CZ)"G@"R;KB_I%;/R> 7P$D/:]O::< <Y+G;M-([*E2\G:*],-P.E<
PQ#F4%_D9A=4PQJ7C3+YTGI<'?11T!B(1WXV?LN4<D,48_T$0C]2J LE@I1<A$KV0
P1.N.5A8R.%*ZV(7$'/X21M4GPIVM]:L'([??ALE(#.=S,7C(HSKG]OM\"?F*3>P[
PW<;M@8S@%K*]D[/OQG3@:BN5(%[K; )5UG-S /W)OAL.NPY[]/6(&2H9$!'P;D T
PP[5%()9,6U@\))#5Q^KE5@?_"T-X+)LC0_'Q9MKRY+]:1II^C)O!1HT!)G9P%#/<
P0HWEAD$P@R;P=<3?2'!D#\IV%@#N JP^9,D-(*\L])P-6@:Q5SFJG6X:?]'(A]*J
PI[W5J!A;!<E4@V6S[3R%H&DWP"$ Q.G9GT&WC* 1 <=>,/X$ACOES*PQX)ZR@-2;
P%D0^H!\5S?M3B$Q:'J9"I0C_[)6E#=HHZUC4[X_1-8E8I^OL7>E7;_ZV(%\:D)L?
PY"> TSUF/5:AC1?/I6<QNCVP,&W!6AN+/@'[3R:AGRNV_W3J1P(/#QHD0688VL7S
P@\*QS<CHR42<(H_R(EOK1L&KV2<03^T4C!Q'9=[%^YH 71;PYX<4T77U+/=78G09
P/3&QS".LA (G>4*0$V5J,S#;(E@0Y8>Q:XR^T)"L8T]/AQ=&Q1$%\JXKK)_<=':4
P'FPP6>_;&<YK*8R]U/I;JOS_BJS^*RH9,)BJ,'IK<5(L>7=D"O9MTDJD]VO>%35:
P\4'(Q @%]'AG?J>EM.Q)IYJ26H+9T;OUZU-B925HG+*9VB\_!^#\1P31A!9 $)%,
PA5Z+.HADO)=B]U13%R3@+6KO63X=<>>JVPK=HVT +3\8@K;VBV/Z+ 'UT@/>1[I3
PB"-&=J;_O!,8:Q5X<3D&/10(/.#J\RWYM+"K%QHQ4;^(N#\YG)8UWF!.;MCAA0A1
PT+CIL"A(M6]]@:@A[EFT?"'#5^AP!R<T[J)KOK<ABM85=T6_YHL?T560%#8$1R;[
P.13NTY5?\<TE S>!N)LDAYD!,C*M*"$@O+8 "L8!P57 $5%(0^'G=W^WR"P#Q>RY
P7)!NMYP3^W4G.\STH&E/=C"B1?Y-%V>0 2,#IQ[3EGUS&ML/$V2)]\T; MS.*_3'
PDHE_C_2.'\0119CG,A!&CMHJ5+"?7N<QD&BIN]WK-Y(ZDRKQ3\OC:ZDQP@KQIF'C
P,U__NV0;<N\^P6BG.GJZMVL$]+GY&@%:"_'0^A;%9*2=:Z36<%3TS('7F$+-H0=L
P.I7^=>XP:/K;H_3//XOKG/)M \7BR-M4TU?\Y[)LI^*$D0#Y[RM 7@9N*GB4FJVS
P<#_QZSM)L;'OOZLW1'Z6BMAQ?ZK]=^H.BD:F-*G*QM/A-C$%$<!!S%,Z7XWU!R#X
PAD1"%SX8!KX!-!1VO/JMD&L5:4<U*/N9QJ1HASCFP5=$)OH!7N?H+3.@]A+X8G3*
PNJ4-I)6TU72'E_R8 J!SZIM+3ZYN KK (ANCV)#78X?5(-=Q/8#P9+/,MI[A"1^$
P9O.&LR?(:]SM AC[";\'&E"?3YQH]M\"3XN;03^KU8S:S:.PH_??PO;YC7@/I0,%
P)68FGC\_S[98;0,_R/SH&YC%Z.L)0*"K%SF"-;&]S]6&VCKK/A-B;8(T78&/2XX6
P1Q(AO4*F5?!S*#@(K8I9)$JG0?EW'KJ014NB-:M8BT=5%]" )?9].JCLDXG>A1%?
PO'E %<4H-DQ'BF0A"FE6_EH3PB5=$3"O",5ZAVA>-@CP K )9FP(2H YSJV&%<*%
PUMJ2I;XF([/HU-@AS7B6,98Y(2HH$W%01KPS(4Q$NFS2I(>%9,'\G4.#FX, 7VV)
P?G?H<4_7UH#R74DKA[J"/WB]TF56^I-Q.;W<H ,C+H5UP5H0<V][]&X(G8&>!.7G
P9-:D)DS$=U@ZU/@C?WHH2"=)H3.!2G0JOPT_I:H=5&]ZP!68L@JQ;&M*30!T#4][
PAV_X'DPH><7$@8900,3YE)E "\JC'Z=FJZE3Y4SM>>8TXMX.?S]%B^1A12SL@/GQ
P/Y7!;T@8Z9(]0CH#^/0<3M$HV!U5?/R28.N0]VL:. W)_J A^L&>+:)68*L/(#(D
P>^V$Q<\/PZSS5L83 <8U"2L95)P@MBMFYU!XL"GX<^DWORA%Q?R70B4J*TGV9-[4
PF)_E/.!7RT_94CZ:FS-+RU,3DQF-4"I'=BO[<<MDE[N$9+/!K ^D3HX)RCHLWQ$8
P2>P0FWVBU=^M&JN*-RB!$P4X;^H_NSF<9YY/*%:B7,!.U;S.$5#B5:8Z)[/7G=>F
P))9//5[O4:F>#Q9=YJ,HOP3@/OC9'_V)SAX[$<J']\B>Y/_]P7N)%?XT"7^7:$%.
P&T)!B<A3]Q&30I6 [L=[(OBG#45Y7;:OS^_'<#6N?/XLTW[!L%5V^*J/:&98S$J0
P,U=<4<%8BKRK$K 8<MSZ@=PY^[_?-+. @P[@$C8?H@S#0*XP(G6S/C'I 8\KN+1&
P(>.'PI#7D%S[:_RK\E?K"SIC>$ASLZ'*X4I?+9[XU=#O9C ?YX_X:-1AM%"'&;;O
PI-S0+ER1[LO4M/#G3C@91#F-#;N2:71$:M=U7TW!\HQQ[@A=$_@K&]$E8VPDKL5S
P(,J4EK'$U&/?4I4Z?NM@CLZ@T>B]X3-SH,)W$/+G,M1A0\26'4%(R2V@P6@?M&6@
PMHQ"X?08_.-07&9UK:M\<S^%ILW66AH%SL&PQHBIX,5+"DZB(]?D+".8KV)V>E''
PO.$0^M<LX#HEK]K*JY\FD!+CRNYDKLH"OABZ?$7WRMA(G=\'(($$N,37?;&1!F?>
PC+_$:00R,C7/JL/KM&IONMZHUB)8/=_@#?(Q"32X6&9=WV7=+OEI*GC9(+IV'B2J
P0BZ6F)YV"L,'RVC);P?R:<+%XTS'VP]>RA%Z;"Q#!\CM\R:WQO?6O]JF7&(R-EZF
PGH2ZR4\X2/6XED/-4(F%Z>X!QV]V)40E2Y)73\J0QSM';<X9_RO8$6RB@S00 H(I
PMN7KJ] 5XS7_?#-C&'%U?PE_RREJQ=-ZEFY&=#3XL\^V#1I'K1KJN[D JH:OH5VA
PU):D6"94Z15'G<!GF/>/;DFS&])\BC+KIO?N#8SA$L0I$<C330];00$Q()DWSXPH
PN32$V1,*7>";#%[\OJ %P2IQPKL"2^'TD/J],A(K"ZN@,C?_0:0->+ ;@+.AE?&O
P%AJX!MU-_+MH&TCW*%ED-O7,0-5QNBUR',!;%H;@DM@WU;LZ9W\-P]E!R9/!O'_6
PU1Y9K7FT]!FXT5M?'B:H5(9S,OA*\/J*2I_:W*(,]_'LK\^:SNS-"]O%QVGH,H**
PDB-;I\8JDOU#7);#.04)1/UV5"7^0N"TFV146@V_W1%NYPY8YK8XL<.*ALP%U=#5
P@BL[,WA"=F=0G:]?.A5Y#Y5CJ:'XMC!N:;B_+6#RRJ/N2::%0P05.EMJKK+RT 5%
PI/..IV.ZJXP!9<00VNAG:5X^DDKKW>'@6\O;L0W>F2)0X&=VC,O 7615BE9ED6;.
P;_X;;M3@ MS5_X#Q'L9(MK%8PP((WMM#3G1&'.*G3>WV#+QK*?,*-92TB'((S3S%
P7";KXS@>J) Y'9IUX'4ZZ?)E@4[J35DGWRC1H73:=9KMU7)5W"-^G>2W%(-J]6UO
PU5N,&UPQG_:^7N;)K8QK[W6!>,@CW!&P\:)D5RVU3WJVE,4&T]5=!:^GE,) RNBI
P7@"BPV51KZYE-EOB[Q@< Z3+VPPL9Y\T_!0;T4G+&!C_/%XE/P,,1V<Q#69)0;\S
P^F7T<OL3V[91C 5]/-TB;1KSY-W-V]H<=AX H='F)4 3 Q#P0UAQC(!XKMHCQSL9
POK2] RS+$36PT>R[\NV"UHNI_N\X ;:V(WU*_T 71Z'-<5(V9!CWV^'W9%";B1RK
P?6:QQZ!K" ,*0"RJK'@V.5G7_&#[FO6DY,$D5MUFANS!C&=]?(AM5>VZKI?5O3KB
PD,>_%,-5ZPC7F#P6P=L;;Y\Z7/G-9T.1D@W+VMME>0G%TO0%?*LX\V)53#T=T,^0
P.NE1]H<0+'^*\*?2G$6;W3AC(W^PJK5L+6A4X95R<7)5VTC7A7R3/;;TA;S+D*;S
P#+'+,[O:QCI@'6U!  K!0EC#8C _<3(A]E;N@?TN Y/O?MR7@(5<X^DGJSV+HU.G
PJUF0CH2JH7/E.W=KXGJ=?^L30_7EA$^F(Y("7M'F @^>",^+=[KZLLMA+P5ZA2=V
PP3EM##Y %JH%D?\70/0*6_A\=1N[QXI?5:1OUM,8;;H1][B<O[=ME)]5+O2X9% \
PP%([CA[EGGQ\OYNU["/L[)X'95,J]U>:]?(M9;D'-[JRH'_[<;I-CWVMS#=#@N Z
P5F*H;=SM7^'@%.*?%CCA-0M"$J]X/Y31W*Y=*-/=/I[NQC13EW#/>Q2UE5VDT]-$
P"SNI=H@X@7E-PM[WYW09+A6)*KP)QRN5V46;TSR"LU\;?$^SF,*?[V6^#IH58RN^
P4X>U\U'H&A%2FJO=Q+AO>NG"K?%1YZ_5 /;EJ&R "02)2BAC.*U(%ZQ8[ESNC58Q
P]%2SG:PA0E7HY&BFKDCOY+[0TRN$A[*3VTC?S)@9:7A67^B);02^FU8&K:'X57LV
PPZLL-OD>0].\&&4KH5QQ"OD5# 1/ X6JCW8PUMKJ7>[YG,3Q4($#F37^97IDDE@Q
P;K ,91+XR5_A49G6"JB_ZN.WID+G5?UCK>?<)S#RVZZ+@3LJ>EZX)@H_M>Q2=$$)
PT>1K98Y/7!GYN!319VP1!50]15YNTN%'NVO/;8WSL8"1 #YMDX;3\5@+W0B'YTXL
PH?2@?)R/^%J^MKD-LNK<7/5>V^KS^H]]4*M'09$BMZ_(?$!DL;GM8QHA0M(:9'S=
PTX,6/Z4CC<\<7OP'Q)KP( CZ?L59\A;ZYX@B/7H_\XAVV^]9:J=FN&#9QJS#^KF]
PA@7'WJO>^.F_&K/R^W(@)LR20J6\.68_8?,2Y/][2F4"(DU="+,GK[_L'O=_;'EY
PFI71?I$# PD$REC:"=DBN,/7=*(\@X2"U1%)K3^<Y:_W@4V;^CSJ\#3Y!B:AZP#N
P1A5;KM23+6V54;CNS=",3^!5=W+"5 ]-5VVS4YKF 2&\E##9N-JK/!F4Y(M;/!8#
P7K8_^H:Z6L7ZIZW&/<:\4@DQE":B>>\;,$F/V4[%$M<Y8,.UG^6<U(\L&U<&\9N 
PW3>+!T\Q@:.(\T HEMJLZT=_5"/973G0 F<8"=]LHW_S32'XJ-RXW%SOGP$+1 A/
PALQ4[P12 *:^'0PAJLQ T.:\QS7B]G5&A[?5[27N>?$6@,EDP2-^KWNC;4NQ 6J_
PH8"IUPRDZ1,9MVP'X^V9<8I3L.X(G94Q(4U"L?L+-=YT_HV%-$!Q!O;>J&83@?BF
P] *"SW2/:E[W1]YI,Y</J2I@6M3S_<UF50PQP7H2U\5G@D=R<ZI$&B IM5#7( W/
P2I8\PJ\R^6E#F;87I3PM$((-"Y&N2<>_Z0@^-; 'TIAVXP'Y3;TV% &M\EK\+I-5
PN]*B(MO@O'EJ3H;.JRFF@-M"M4>\FCL8N<2UKW4IE=MX7A!K8<Y12$[8,?E>0:ZM
P;EG_^1?SX&.@CN0C12 V\YPUFAB6-Z5TP4J".#+U0_LGXE> Q![J]>1-F*0!5UIC
PG_7!L@Z*+&:,4BXS9EGU>Z^;D*-$%<4T*I_?X_@TO97/$?#,.6:X;)V5YAOS,8#S
P>V>E^WW_$O6"67HBLO"G>/FLIP;7>]*GM[Z5[,6)TYY#-BDQH-:2;D8--[YM5E"@
P!)VLMG$^T2FEA@8WC>^AAU*_#9Q"?3SH)!N)7_O [RF![9#*W ]HDA5M4**RN$W\
P;1/$@OM7H+4K%TA/Q)<X"#0V.>T1@F'IED#\L!8L2!RQP@NS:"(XV@974W)%%O)W
P-XUZ@UVL@5D@-3EQ+HI4K6%/'J:NNAKTYN<5OFZ9)M&TOH16:E%-;17K5ZPAMJD+
P40$03A!_L;0,(WL^*9D*2R+%/WH<W\4< '9]4IFD7)_V-T,B>?_DAN@AWH>Q%S<K
P4!%MRP%.1\9>G :Q>U?"0MO6VLN)T,1!BP-F9F5Q4,R05%USB&,5"T:7IVX/=L&N
P36/,&X:P91J:@8L?AR2)B5L>*53C# Q>Z'N8DTD$];\"'RC)Q&*OJLI!^G/7Z"=G
P-LBC"&M,/ +0VHR I&>HY1>D1<98&3M*T_PE_ F&"A!:4.O5/D?MT- THU-)EJ@W
PC1E)\-YR&\-KQ#!&D3MM9RF=[U4&-BGX'/B)Z!?4?7:VL;E'Z' 2*?,&R9'O&[4A
P=YZR]DIW_J"*B?3YD8G;_]R(TL(X?I4')TQ5) /<V0 YM[S%^X3JKVVN.UAEBN:L
P^=[MJ67K;Y-@,5'-)HBKK)3E$W=%+$$61V!Z?5,WN Z-<W>&A/UW*^Z4"V4L/9*B
P< 0 VL>.SQFA)<^55*Q/*[%8B&#(!9$UNBIK$L30H:PE>$_!]MO<,=O&XE&X&WTG
PJJG%<RU_)J;JU>+YC9BW@2]C"?7BR-,&J*+$4DQS,"8R2"%UHO^WRTTH!I+L 1\F
POT>0_B9PJNCHD ]W7G7#<U[*DPTV,]-7B'EA]#@JL?8'2:S QBBB#'XB]*&LFXT4
P7+LK M+5WZ=&Q&XE1=O<L6R9$U/N,G*41H.O1P:L7=KFQ(E:?V0XJDQ71^+M8(0<
PXN5Z@S1 U/P@;:, ND.(O1R_NSMXO]PB6V8+)OLZO"I7BU>--WO@R]Z?U$1/JSBJ
P8E2ZG7?#G3E_F$$(F1@DMJ[%YBUO8N9A<P 83U>)WA"L'=8Y*J>/-3+)&+]_5 +E
PWSGIE52.Y30]P8*C&Q\@FR6V9#&*YVWG1D*9/B)5K@%OYGB7H(Q.N5T#^QN=1TFB
P?[-(?5!^KC#2H3M9\GMO"IE;#H4C:SRMFLCR5U-I;ILU8 5SB%ZXXW+58"5ZX0P[
P.S+T<4UR'"G)X=JXBPS1)I;%%2Y'&0S;4$>&K-9Q(VVN1!G-GMN/52321NP(]X,/
PC4KR34I=.RXU;A,?],".S86'Q]W+6SF]2:&<9)=Y+5#Q;N=I:W_OU/_QK:0)^UG>
P(9JBNC]>5XYB)7(6JN?H\(O_?.E&V(RKH50$C^[$P=9AFP[$MTAR24C0(D:NW(0+
P^V6-[>+4;> <(FIZ239"$CZP=B.0,!Q,%M_K FDZ//X#;]X<KHV>9B/T0%R[8RHR
PQ5O_MN2&7::WO;7#D))D7%!#[P/^[G@7FW-ED[N<S:>J>&V2)5)BOA)S9\)K6@':
P^9+M!G9U*/_X"E74#TB8HOOE]6Y(X:98H?1(# DY;[*R]CG'I^RI6DH0<*6O+R"A
P/%%5U-MJG5#">#\$M$P^GPEQG:S)GS6AHM+H[E%-N[R&8?JCQF"-_9ZT3%$]^J.?
PT8LI)1#)_#AUWAXX1*09;'>%JQ8[7V,)ENQ\GABM^Q,Y)U]1"=2M;UK2[75,B5V"
P@-7IHCA<>?XTC;EL:JM)&E _@P9_.D8)$J%0[$_"+YSE]!K#_J!J/8_IXE<0DI08
P$L8^DM2%(1*_!*W:Z7G^&L7?P8G!+].HF(!6MD#JP_UUT*%1O35[T*'IWB104@%?
PM\1DXC89;H583-33F52&A#@4TPH#^4,;FWS?7H"F+UTE-MI^1"X 80"NP&R)I8 B
PA[&5QM]4\&:^KW'#B35'GXL@14/MC<"+]'Z>V T"78"H/*<8@G?W3%MX)S>0"YN>
P@/L4^0>!>6P.J%K5=\[D[3@7@P1]IP,JORQF3Z<Q+"%.TT":#.NVW ,#'6",VRZ,
P ]4,,B$.KTY2[;IKP101$ F^+B][ 95/Y)V3N!M*/M?=O.T^1X990L'UI%=L9R)E
P^)V9S&*+!-TGF!T=^AM0IQR&<@7C,6R$6V_.XSAN0CA'49XE8+AKBI5[,6R_&7*0
P.,>@+TYH*DC9YCP5(SF&U$G; TYXJXDKR+MK,6)8D$??:E>YF0[9AHJ#<_N(*WBG
P1 T!L/:J/]:*6%L+ETNQTB@+8TF>KE-K1FY@36DN,+DAK$7,8C;202C0OT1T[L=4
P2F'H;,5#D4=5(IYLIG<$* I?%QZ.3(<!AVTB_^RCJX;-_"$7GIU5V6\%49";L$&F
PN-'PS_/MFQU^=.1 /(,NJPDB$'WLY\K5I/H&6D70B/2(%]F*QB12=QD;$[?WQZE9
P#E/_&Q8AZVU7+$ZQ5*54_E6+JI:9D?)Q^1Y? U-X+VXY.3/Y$Y2ZSJ;NTO=PE0Q.
PX!0;S>;&_Q\O#-U)&=&6XJ,0L4Y/OWK9= %[*Q=/B%=0['.3LE9K4[E&+R#N%6'N
P^ E^5@HBQPM&)FV<TO"Z59"+@0^9!FZYJ-:0CM0I0,\[\X\.Z_YLA4#>62P>2O8)
`endprotected128

