// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// File: uvm_dpi_helper_base.svh

`protected128
P]0: 5! I(A&F&"X@4#CM2XY4;;IHF.I[+: #JU2!*I&["-"Y4#.Q9QP@_)[^MGG#
PMV!XG\Z<)'QHW:Q]V$766RLH[NY3N4%KCE+&3?&*Y!1CH?37;$+[*,94UR=C!%&3
P%Q1Z+46XU7,!%'A[ZM"A!ZT\@XH&PN@<W:S5,^S-6O1"S9J]HTP=P=Q[CB6I^;+:
PPXGEI0D?YD5D55W&DH;A][)]H-3ZR],U=?\(+P1C8!#;3J(^4;S4QF&,'XDDWN])
P.RL[Y >0<V1X, Z!(:F5--I7]N1]"5Q\]0$&E7N(2NP=!S4T8V%B83;,%?Z84JK+
P8NM:T-EU< J;U)SL]1LAC#6@?F6I,4^@60/J\>M^NM+M)0>>:-1!)90!BWJK %-3
P&RP%837>:%!H_3Z$$Q&U">^/"V *4F*2&&X;V3+7[MDC+)I3U@WY?<LS)%$$\$:H
PHM(JQ& F=KJL9/]-#B.IM 8M4TT.S$-A*LT)*VU4^=FBH[.YP;_*/KU>>J'#<2<U
PTJ7.9LEO;"=KC%<B5]GKADC-+L?_?&B1@QD3"+"649IY9/AU.7#;6:,.RHPY^O)&
PV1RHLHIP^S,YY"O)/+'U'\6$Q_NSM,JIR8SEX+AOH2>9#2O0LC_Y--PX B_5/Q_>
PJ;Y():85\ 2X4 \0?R0)D%>_,W%C^L^"'0:=W0HG$2>G6T2*+6E96'E*'IN$DD9V
P 9\-M9_(2_9X37K]PBWOY)-'HDLU%!U/N8GVDMX*R94P <,X5$Y#=0 YHD?1:RC0
P7##N2>QU\"Z*X,KA7*2CD$X;F1*=5\J:M;=V*1C4S"N;25>@JH3KO1JJ\>DT5Z*2
P,6IZ>U#&"C0NP?9KGKB12$&B=X$4&563-U1.GYM863)($C>1-)]1Z'3+A,9E;G&<
P>BD@YB3AH_9_(Q'&PN>?C&%84X5L:>/R36E_/ON+D-2Q$ &.(L]INE.=G?]19FM=
P'SO$V6CE1.U2Q.-P%8%5^[_!7('WD28ZU+TBWR8(#)T,9=)YJ=5VEC.[XJ0'"/V&
P4HYR=]K$Y?V<]-H.J*ZEQ^JXK+)SD[(4(I'Q2\\[3W\%>%1\_GUTCB$UU5:?B/"<
PF3@#"8F@#L_# /,B?XKRG+@V4A[.^ %MFQ-FA[:[N\+N:!7MOA0914?93<+;-),<
PYK>DW)+2/*6J^OPN)(X52R_-<*793BS\>?V&*V_I\XZRR='5W>&W?&!R9EG@'ENE
PG.+]Y^D[ \O-Z2&I8G&2]F3T \A%-Z&04K8J'RL$ID>UV@VRJ&F\^HS+!L?M]VFO
P6R>]2M@Z;'@%)KMVNIVWKM^X>]32U\ P:#=#"#J5S\A&CTZS#MSK4]R[HDE1<<AW
PH-O-:;,"ACG:&=55'O:,YKG?RS$H*L?3PUSOA7'72]%95)!V3]+M0RHY]52;GQ'+
P93[0G^'.E!>W:82R#/&T,R\ZYX4:OARV.6[%VHV.>6,!#P!R_\E4QMP-%)MKF=B1
PR['691MA;N8RQZ8%<_=A@@W1>A5W;MK<]-8!AB4[$!7U$#K(+YPEVJI:W<J3WIN[
P)S404(2S<AURW'2PPH;4Q41A)DFVV/Z>-OWS[$3C0MG3V.^(B+:,XH#RT?CNOMS4
P4KDXS@1ON$5 ,0#9[Y9\9 3'MC=^5V+XR"<TAZL!*?IO56+7".C.@NR,GCF4+19T
P1FX*>,:@O=6N&@6H@R*U1B2WL^!(X>/:T^30/!@LTZZX4O">VR#,Y!65^%6.803(
PF+$ 9*A1!^I7$2I ];4Q+A$7'H#5PO,.QC_.8-LW,SRRW,Z<JE.,!#WB::'84C8!
P;HZ(ZT< ><J*:6+!@4E/.""NOI14_!^#]20[&).(CH&&$(?;D_I/+G+N0Z)"?AG4
P"V@/A$(9 ):@/H&$G4@7[ 6L/"N$7T,WL?:GIN:E6A2'<OC^.%K\A'%=9S-T$^+;
P:FVR,)3T%#N>['WH7;S**^Z<]!& U?_5=YH2P&VV7;&6?*U7@#P=J3?E+0[#N,0A
P<6/@='B,N64BX:;H&Q%?(8F-94&0@#9%@ C8@JASLZ%V7]1!G;;#A!70W@)?=F'(
PS0A.U?8YTXY.)M%-.3B2@XQ_P,%/EA_^*4E1QQ+3^^W2[Q*5;&P.2>P7HLSF!:([
P,V#\@\V\P;_K\3BICKR3)YK[;HB3 "SV*<LJZ_:\2;W&>T'.2D4#V!D1YGNGZ>;W
PMX#Z!@X+/]D6B'H:1 X+R5=NR(5U?98=@.-TK\P)W=A-[VQR]NP6\K)P6JJ4!!@(
P]T  \>NE)RE1%28-I1CI&Y'4,@^"?Q:-E [H*?52KGV+_&QZ'&JK@P]@> X_;G$@
P(V.\J9ET4#0>Z4['/-_'Y.=]T*!;'324^#9B<'QWHWPC4ESTE&+4=24B*OZWT.YI
P+>@HSW3'*Y02?<)'/8@]2;?>*(+U0-9!S)*":^1 : B>SF(C,%O"J<09">2ZL91=
PB*>FXB! /-2$&)N1ZKZZ^=;UG"LS'ND'Z%N)<U?V:\274NVA*-%N+C?R#Y'XLBM#
P$YVWN8C@2SL06GL;)!DEOH2]9 24H"]NU4?L $CF@*^;+Q-=_-;,G?%!OA7Z&GBV
PAM-X\1GM!TLIB!S]'131JY,>5)OX>=\4N&/F8 '1QE?2A6G+8GC@HGM_0U8843K7
PUT1J>\:JVB5K<&">P#CRVHI#MV] FU2(D=WL#K[^$>T[S<<+4X<EJ!? ZT3!*K*!
PLLOPU-Z?RKU^R#F@4D%0?CQ(@SM&Z>:E*&HEQ<7Q0M<QM8A%61<&/]8*Q52)7FI?
PUXH54T"W+*<FY?JDD7*@F6HR*6:&EB!*ZGNI1OQ7?0T&O6GJV,J7&QL]8I+AN/!^
P5P5779_(4S/!17JT<BB78]?\\'F"[VS @TTC9K;2[]F^.!]YUI>Y [*_;UCT5P69
P%FK@89H15+<-C[M&<"3Q;WWB74Y2>#=;%(0=EL&*;A5T<HF1Y=4Y&;31X;X]X%-Z
P%DQ1F5Z6MYJTV%9SGJX7WTLUIU!N.ZK6_]T8D><JJZ@&/HCFP5R=KB!74EP76UUV
P'?<6#.@C49T/_,GM=I/PK16O&#W?\G_ M.6&91P)D0E;L X)":R<Y+*QDIFH>QP1
PB9I: $;!2:D7!J\REJU27 ,)8VV0W\2U"1;9_/]V4D=;CBE7P?+D6/_K(Y[1Y(JY
PAR,& ]]>8RV%V=3!:)8QO_.ZCV755/F$+SXH>^BK/OA1>%?J'Y%)!D:4@NXO:#5-
P3@;2QNU!!H,N'R.D0$NHAVN.K\6<!"FP:WZ^?^KZ_,HOE#I;G$WV:>+4!HW6SV0]
PSRG0BY=2P&6H[C<$2E</'\8<S!I@#(.YMK][IQ^8L CX'2?N4J_,L2=M.5UB)-9;
P!FX.]#%!9W'/%V@;4IE:2S N^@:['_-PP&(677"T)?*^:0;!714L.RTP &*58=YW
P_*]V>)''O2/\K2;MLYH>Q&R.1?QYN=67L/,@LX1VQ1[5JP(.I8QM-K['O?0(O".?
PK':^*JY#U31'UL&D:AU>4;9\ML5XJ',%XS-T%3NUL/O<TK<8.EKZZZ(JJCQ=L^39
PB>K?BBQ+Z^2,IQI/$=>K9_[  >7H!XBMIBGKV<)4+1B:7Q)$K)$XP1%94"#>U,!P
PE\><C%=!W'+3J6(OY%$9DT]G DH5&:;"(0_F]^!2V5CF+GTI_3H6.A&5TYWHWFI*
P5^2_NN[(] ,=WBV/(2UPHV/P:B?WA%-=C*AW2\$>3G$+K4LUL%$^4JA?=W62[A(O
P=RN/9CZCAIV>>Z1D38>]3XA2H3^)#*@L0.++_G[=N FS*JM(=NG*_=O#\)]KLS^U
P(H![Z#CS%+7&F^5_K: 69V[HV=I=2&#-XF6QD'T?K)O".U[]HTCKT-FCQN27W5'D
P?ISZ.^AHP)L2S45WG$D68#'WY29RN@?5RAZ,6]:=06.0[PB?7RC'2O\$C42 .V@(
PZ_^Q=C1J%R)ZT5R7 ,[];_.VH7N[_1U>\V,O1R!.UNE"^:9,?=<(CF!&HNKX>4[Q
P['A*UA9H\5T+AA*/-8,F50O29B$Q5SHSKD]Q$XD# :?=*2!Q#3O]*8F7M^RLH>U5
PD.0/:)%CE;_##9%=<]IAN1(^$M 32CW1QT' (_"RTEA$,VJ]T9*A %\9XAOL*Y_-
POH.KQ-IS(Z&A*MZ>.XO964'F6P8.(#%6,4]#POZ?8W=>A>3$2I"+!6P@?)I30"//
P[JRT!,_5@^0+IN_35'_F9VL]W[^MN,/U8&Q.)=+4'U?YT%AZ PI)32^AH-L@#QE"
P&&&P7\!_1$Q!21S\N"8CRUX1] :H !XS^EB6B2IENN  (0H5L?BY;9PWM[5!>-O=
PW6M1+V:]9-,^?^I(7'FY'R*C4"1EC2\90WL*&C^7J\'MS#,M^1GR4WR(D^N*(JYO
PRM':.FS!F=(YNW2+4!/;(@6<1#?+=16_F%N6EP3TY?G46X!9,.X7-]GOO>2:R\_.
P+"D%6G 6 )!$8%5M4_8=)L-/WB=)@FZ>\A6=%\!&U5WB] .KT[#6_X2+FBM2]<HO
PT(^ \/@.>C3()^X]"3>?FE;*-NL8N]DHJ5-YP+\!8Y3/9H>JJ53/^-D-]CE.;V)D
PP/1E C;5QH"[ LYG==15O%L1P,'W 2@^%[ D^?9"#U"I/:;-/3U0@X2,=<]^5)'W
P<1WR.0'(A$)Q [&",SLFE@,L684R9WBP_UJ H5Z2ZA&&4?99969<$Q'[+@6OMTV"
P:JB@.+C=-&'O)W>_G[CH3]+$?HF5F7J(N J%8N).+V!>V+@>G!V.#7/9%#$]4*NJ
PSHA.@EU-B;[1(_T?VQAET<8*3*NPI?9I/>80I>-NIC-G)V3"^4!=W=!AMA^*!2!U
P&PIV;6%=H^9:/.@66XHS:95Y%O?K1WC#-:VP$A4BEBA*#0ZH$]?S-/.OGOIIVUY:
P[0#-PLHV%4"HU:LD)5.2H;!_PE)@QBYDQ)VTWUJ*Q%B;!^?!)ME<!72_RU6;*\GT
P=?6=P:0)GX$U6;M-9^*"Y"<"(##(Z+B5RB'4:FZK]_6.4R-8O^O9W_O_;I&PY5+4
P >ZW"C&8ZQVK:0]ZI#>A^:<F02$$^+YZR+X!D2+#V%Y*0F"47[_UF#@Q7?MTX+AQ
P"V%$N'C;P@/)\DO#H&I\)(V#4(V/:!#BG5MSCOT^6XO.,D$\029;*"^1^6O>V1-0
P1--Q>3QK[[K895L5],7$HTK$7]JR!BB4R(@*<PC8I[/WY"M=YNZX+7NL>+8U&CP8
P/U:C01\++.UA'O(BK ]D)C?_M.@K2@!,F?CA>6^<^[FQ)9K Z;>;N;#?S[U48,M#
PQM_:O^V\_<3X S*^OOJ1+WDM#8JY^$PI4T*H3^IK:Y3/TB<6CCB2/^K8JV%2^(/$
P^%-BFH/<[3N:/^#%28[7OJ^:9G/K 2"4T5TH>W6]"W.P$YW'E&EX]TDHKMYT+D%[
PW8VN62H(^8"VBN%0?ZW-L3_:7[3<% 79!=1\BE\T]TA;\@\70@%" ;^^NR9YSEYN
P:4"J1)B3=E-IP6#/21U;1L^ >6+&*+RIY)$H_"HDGML.KN;(N*AIQ\C:T\,?TGSJ
P9VE.5Z3=K+&_CXV3O]GIC#AC*N:G$N()R> 0;+2'TTW>X:Y]^7-]H7C]C,NH(Q@H
P^@[-GP18'BW?"<28I0 T[\5VI=3UOC^EAW#!!?%V^5(RN*;\+.9M-*^/VSG_.G&G
PNEH7^SD6R/W[.KX@8O-<\.0A#27$+G&@";_6=;UY-12;]F;,#C!.KI-TKYQH65 T
PQD#%MF"E'$D Z'+V7&V'_+<QVDO_I+?TC65G@PO&F79_BLHN#5;-'Q#8[@8 YR<8
PL+YV9+(*70]0?.;JO!5(@6W0Q6SNR4>TI?VFV,W,2+3^@AL89.]$><V6#>.<HZ^-
PV=@V/NRCK<&?CULH%[WG4907VKM6[3\[AD_$M!UAFU;6IC7MU)8SS#YTL="_M\O=
P]_W$4KZ\N@RP%/-J?2-TBP4:&%BG<[LH_"8R#C,$(?5,@T]:,++GG\>_9'?I(;(T
P$-<W!#$<<G>W56S -K!(.=1(\G,(MX]GV#U@->1_J0):/$$WH&7:GL_W>UQR $JP
P)J?!P #*.$8=[LF>B\V@CU)8QP2V)-I#:;CCMD)T-@TU#U^>TN2HWI- QUCS*:AM
PSC.]V%^F#"/R*%PO9NAXQA;Y(>S8/CG>-$'X*'F;5KB@Q80, ;VVOMJU@0^<++(P
PR@)-*"DD0\.>IT-2UP3R]QQ_PAF]@<-7BXQH9SW#X5/[>"!\57]PO"!!K5XN!*7T
P22J3V%8\]9## #ZE3$7%AR(!RSL+@U&K(Y(^UN=XZU)^J?\_E<Z""?TF+@[[6*;H
PM9D],F_++YQ0)L3"9H1\X.AXISU59J-M5*:[A"=H15Q@$@%L^BM$SCD 5_QBS!/8
P71>&*_;C5H*!-==5WEB&F0MDB8U')P!M::\(#SI!Z#"8+@0>,265_QN5%%3OR1/%
P5EI?N@+*/?.%'TE"PF2)1/C\'1KE"(-_W)CZR>:#4+ $)":N,*.,'UG@*=>)JQU(
P98/PT'#\ XJ+(ET; #:U+]/F6A-S]2J'BZQ2QN+X&7^OJ@\5B'FA31+B&%VQ?WS4
PUNC2[G>#VJ9AYFUNC&9=')1-TX]BG5Z]B)%Z/\W3C-<^]?9)*WZ2@0OE8MFE)6I_
PANWSJNS\[*YDS?'U#UN#B O/(Z ]RK%!76!Q7&&'X7V]N7RZ=MFZ$T8> W+Y^\PD
PV1/_&'%C?OY1F<RFOC)#XVR_ZQG&Z=*[OR-,(N,=):L$\SE]@=_N^E=KRI>I2HBV
PH>DWGA]1RJ&\I=3^N">P>NNW[8FZ0@TS%0U*NC[EX]-@[X43Q_"-MX9\9F]WX77;
PF9Q^,W5)>51URC)9A=BO4H!N#<)OS)5086.8B_^AZ]-:L:52NY\(C3</0E/A*!!P
P5!!0"S#4$O4E=^\F7XP4!(Q'3"*5%"SH&IOMBVIP4^GXR^6?QT;\TR[05BG;=!B[
PJ,VD'RS#9QOU8,5^N9.^:THYHN)W1/PH^]U2423RHH"F0G,!O,Y2=S.V6:/5,0^#
P<J#I5_';3,Q=5U['@5?#K=KA'FA78S(Y6+WK;N,UJW]B[XA@(KC?P%;SG+!RI@#(
P7N;VDNZL'@NH'%# ;QHS"XKMJ\#\UVO/\)XC<=WWW+6M)DCG1T"[U&B!['^SR0*.
P;*VA9Q49ZSVK?Z'!PU_Y $Q9VN>C%] %4M*MEZY2++:W%M;^%HX-P\X*1(@ !A Q
P,T<R:< 8RY7WH?W]IIX((?>_[EYX>;&.,N([G@](@T46@ENK!YK#T#=/,%UKXA#[
P]F)%JL)INFE8<X434?HS3_T'8A(F!Y53U&R3E;V G'-#R#TYZRF3D8EXH.V\6\HA
PC,PY/-JZR#^G"*!("+R;]G.OC4]H)&U;^\O4/\69HL6YDNTJU+N52OB%O3BB?)FM
P@_4I%K<:7<04H?S_:0J'9GDJI-&R[3'S1?.V&XU\)!\93)Q(!(HF*2$R61;7$\9M
PEG/*I1D+BF;"8J#W+^BDNC#GI]/;94[0N!8HGV^P+7&E@4*3A)+0K>A,_W1Z0%7A
PZYFNQ[%]HFPF?FOZWRT!5T1)+R0!48JOQEJXP=SAH8;W:2.M0J;ZD(-FF-?Q0LR;
P<>S\V!M*G Q#?5*OA['#5)F% OFQG=(L AL#!D3IVS .A 'G*X*1Z+KTKD/V?%$*
P3_G4FC5Q/O]] =PCU7B;@69S)LWX"RJ7(2BV@FIR;9<@*EXH:99U08!Y)&@?*7[.
P5$6(&+1ANIM1+WYEW#QH*$DS">?,MXSV;4^,J+6A[/P-YMNGQ!NRAR4#K@":9@Y-
P.HK^/C?,Y8<?N7O#_T>*='/-C86A5MZU[]D27E)5]VO,#J (HN'G-_X*][X_<.1/
P,S13'MF;.QU]HHVAM?]Y2VC7YZXHFNW6QUC^V\-=F2M7JXYT]<CTC#JDD7+*CX'P
P\\-O+T!@2=<)@&BQ8R:[C\QT@FUZMD@V?[@)MU;V=%)[CBPAF[63V=)0Q(?CLV I
PRI0W138>=BC"S!H"')1.J.+^Z7/KPZ*E)4 _/?['FV:2=VU$<SB20&=0 ^&;-I^,
P.*)>4)C@\,!VI%C.4Z[-;P5DUS6;S2\<S1;1/7,^I4'R3D%6Y2_:2*^DNDO-":LD
P4;GMX+);[.,<UBC?$J$8:CO]4P69E^EP-R>7O\ZUT\JX.T_-%WW,0:CWIF?IJ(\P
P$9JFY< S?3KK*=&]]%R!Y]V!EI=X=&0O#7 25_N()&:#WB+6J[,U1XN#WFJ0<\ 4
PN/UC*51]%@ULT_!C?&&9?E S7UD[5A;D+HBJ+^G<Y9=F>,62'<P\B=LG5-RU8Z[C
P?!1GY'FC]V8-:'('$E@!N$'WQHA;Z-TL%@&1W_J=J%A#WTV=9G 0R7V>0&NZ6>X%
P^Y_\4.=BZQP;]3"TF UBK2"/7Y2TGEN1ZRPE@30:19Z@$I3#02IC99F:(5'%D'P=
PQY(@$QT_9>Y&Z*,N!GB6BR=\,3M#B 2=<-W$:EA*.=\'1+H$RW,=CGGNX6OTJJQI
P78VJWTUU/1VY.=A^BFWU_)C.A4#YT.")X:)U6_%^/.S0R@D:_ACGFECL9DS(A?QS
PLZUQ54:*?@!D8]D"UAR8"P6AR&CI_KN2#4;Z<OL0FU1/6&!(GG"!'X%+6O@^#](L
PP7]EC4[1A%YIT0@/A$6M=P553915&M+L MQP!9H!F\2\Q D9XRKHM?*OLFQ#E]2A
P/(8-2IX./S00?L^TC%*DYFP>?T_D2T$[_X<CV/G3A-M%5>]7.7 K[D4'K)GV8[9N
P]214_Y>#6Z<?N5D(/H>\8MVGV./X43<UQ%HE^Z+P=]["7Z2Y:S8T)@:XV!//.N*T
PYTF$"5WEE^R"RGO5@/=?++KU-0N2 &4>]28U9[UAGOC KK#/\*X-Q>32T\X)XL^O
P?J('1>_UE%_NQ<P5!Z>99_/\5';N508V1I&_I>ASG'[0%C19([.>W^>:A/@^AILL
PYK#'#*"G.GO@[EM5*.\XO;+NMBW"@0JA\J,Z$U00PG(0/"'ZNQ;0F7L8SK:K5X=6
P//=LJ-'<;F*E%&K[!XC^GQ,=J]^U]S?<F%/O@XCI0?O1&?W"A?52DZ)6<2HFWRGQ
P7^ULX0#3(+;S)4"@OM@7_96@_-@M_'C<*47D"11_^/V6?WH5Q)U4Q;&\O,Q.OG](
P=%W?@Y?:?^IJ5NNSO4LNDZ> YQQ)/G8KB(?F.V4/),PKE".=C'%YO;GF^W5S5Z2-
PCA%190(%-GS-BG6<Y_5H4LX8,$WRJ&R<WU/K>![F.1ZSI26+&@P=.].0PL;;0KJV
P0D4N1]+ G+$'5QE_"U%2?>C1#"X(N,WZ\WE$M9VT/;**,AAF8>#UL_U&^ZK!C6N\
P":LTSAA:)I[2>X7:H0,QQ:YLQTF=IZ\T"V#H?)2%,T-9C@,^XRL%!;8=IQ[\C7AS
P@_"113">LQ1<A0Z%)XDRF/[(,1>D%]8+S'3^9.PF)<L&"GVA2$"E4(78Z<XDI*KC
P:\P_J'J\!K]"AS?]J#O%IF%EYM U?2,V>C%CH]0"2',*X*OM%^"#KM:(VG:)I#?$
PR5#HJ#+"E,@@7['F8QS=JX"!Z@P!/5:O-ICL0P0!_QM^&W0%V;?TN\)X3'HNK02%
P1.KCG/BS1(5AV(5<(\2_H%!C+4\!IO/"D4%X0G3XP)0G2^'2+A);[/YP>\& 9NG;
P!#SB_+?^,5//+;5.U=9$ZZ2G>^$KM:Z:UV/NXFEA8[+)Z2Y>@QW&YVQPI4/MT<&)
P*%-38G?L((#@1MB&K.D<G8)%4J&W]F)V2"J-S.)WW^02^R]+Q$J.YDA+S^*G*:E0
PG\_G(Z91J.?&Q.(Y5'MH$75K(0*-HLCA1CWQ@MK,;YHRA+D]/>O%_U)W,\Y]<1HJ
P8DP-F6LL+'FC-]5SJTTW/(JO+BT\<1Q!7#B?6Z%4"JRJZ@1JXS9K55*I!=].OS/<
P[T.L<Y.!+IN;S:HU@:SXX0GF,E(L#R5@U-)U@(@_;/,2*R=AR0S,[SR8T9>=$W6E
PI.2P[D=V0J$9QS2&SLW"JH/'P7B'O>[#H,S][/5D!ZM:6X/NT=)U3W+>2)Y9O'NL
P3>A*)=])!O]5*<^EG'EOL4($^F&SZK6J(AZ3M)G>.RYXO2SU;3DL_FR9E.=A+.50
P2# L ,"W2FU-NR7S6M= )Q&!C=M;4%L?FP2ZX]VW]UM5C$MRQBL71Z66WH6IV?\@
P@V]X2B90;'GPF+4)Y.\I+E?28@FQ"?YG'@>TIX%SD]MCLSWTB*$$T4)\(170)\M.
PS@.376-?3927W_.VEWI5+S*P#&L">K1$)TAQ<<&C-H\% U0H&U@W8T\9]@&%+=PO
P6GK9"W\K8YZZ4"9:"(T*AX 6Z;[*WGDEA>RV;7(8O]K^["4C)G]!L6%T!K!$1P)F
P$1;>ZJ:UU .B:L^!8GGO)6CQ%G@>P96X%V7,@:6=7$<&I5PRP?QR9ER#ZV*!S1EQ
P_5BTMA/*W$5QUN8SU/HA7K"&D=%M;G(]N(3=.Z]3T0);8\7YU+(_+^F6=PG56W?8
P=KRMOGSZ<$"86V6;Q5?6@+B;"Y/4-,FRA(K+ZT$J8!LTK[G#0F&B ?Z!/<=@6O:M
P]Y%*^89DD#7A7T\\P@_ZD%9O(.V) FA>+L8IW<4?)O#9GDDNKS&5\L$ZMY9[3'M4
PTN*&*WVKN<1Y@B'B?EFT5G=52NH44UF2 EYL+#6J:#A6X(>9,L"$27QP[#HU(^$>
PNU1QQ&>(O-CACDOIPZ$^(I%%L("3[.'=?$EQC(>T9XM<=MUK;CP,)S'-36Z9#MHK
P 0#X,A\_D+,G>4"7_U6(?]'AG24JDU 0;F,G(6UX$;A^M)YOYD!ZVX\RZ8WYU63[
PM=&HT>0_'HEB$*E[M,SK\/B61J@6M);*XGH(B*]*9Z&!VS")$X$-().#S#&PMXQA
P+=Q<@ 1?1B[5>?_Q$=,80V /YL47S5S:==J#A]R=CZ\1"8F8N77YT\.[AX+VD9+6
P\T5/.*+55ZZ2/!L+!9_P9P=P\3\>Q#Z,X9_1U#M0X$9N_#2BM>RK]/7#/Z:O'+/$
P<L!BC#=SP<@[8\%[/56W\9*DWER?DF]?7./V%UI,8D#".LCFQA=[>1=(B GG6#L0
P!A7OZ8I+;>@.YJ7)I[1*!K DI<LS1_@2-VU=R(\\X03J"ZS8.%*&0+)K>F) 1&]3
PT,'QQ)QESH$FP!*J,:9N0ZX^%%(WT=.JQ7IK.]-47I1&J-FE*,,\@HPF5^J?A9^N
PF<KJYV%YZ)A'63',KN" *X-E[I3=Z@MA1N9%"NZV^6Y^1:+]AKK(W=>]26 BQ@K 
PM^9 ]-IUNQEPOL;]BW B ^?&FXVAM#GG<K.)4JUP3P<;A3B(=(UIE47>AW;,T \0
PV^=A.OX;%%)>N?^#AG9("U4X 9)SO5$V*[WB+&<XTW_>XR5J&?N3IE$EW:B%700R
PN&:/%M#M)AO"HW&MX=N[LVD=8KQ>F5^%>=Z8M8U%&(PMC8O42BPDXH.6H1A3(Z+K
P@B94GW>:2BLA(GK6#2K(+[T8=Z>C XE)";+<["AT3LP=[ZEC%;Q'K(,$&/N1,=*5
P$E+KUY,3Y]@4*$7[S/EK_:VT.K0B6I91'WN2\(!KSGQZNRUA+,]8AJ$Z5B\78JN%
P/^%.H%N]WQ0\X\H5OI[,N]_FW@\^*C6-^.#Z."FR(<2)(+6K/^/V-091JSU66M*=
PXCI*?1KI;WTA[ F@9W2.1" 43Q'#RV'[A1.19RNR7WQXU^I/UG,<5/>378OYK?UG
P800L[GIEEWA1.2-,8X^#J8;%&DB9O!A0X/XD(Z*(/K@'5H0>O8KV7I[*?=/A2_9=
PR-P$[IC^06Q6AA,XGC51>:#_YM$O.8U-5;J_&X\WOOTB&B^A___-8XD<[L-"O,4Z
P$8[#P[1E%?O(02W\U$]^KC[)NIGPP=+Z %5S4<^QP<'/O1BRE+Z38C*M#II:5T[*
P#"8<JJE_MK! 9('K_C93,P[72JA9?LV[R5:>4N@:MI$PA)/M7!RWBD357R*P$OG,
P1[!W3F\<;@)CA)$:&275_,J4;,/Q=/SX15.Y/4JU_WW0<*(X;^KTKD;)E-HBWL3X
P'W5H+T'=).4P@<OF+1<4XI1^%:+N1EG6V$_C9_!GQI%<L_@:C!P*V&,&WIFH_W\5
PH>S3KG')60BDI6/UQ(D]6*3KT,%KJ\7OF3K]H*SZ%?^R'A^B17+H-+3L<4<Y_)Z$
P %\@KHPE$,'7.VF\Q[CLH5S'T-#?U?O!8_IB>)TD=4 K7UG6BI]?M"29$C-O%0)O
PK.3I-!.36=M?WXQ\0&(IR(TGBJ,!.C[.USC<7XXX";\0?@D@JM8KA<*R4LGS>7AI
PJ$Q\RI&LH_TT1!:?RM,W36(Z'XK:^)-I'*UV?&EQ[>]+/](OE%B7-WXO5Q:<FU(C
P.D8N,Q.05EBJ\SME>X0MQC#<_D<O\2-S$CF19I\.?L99M;4>%<@-V[?P;)6PX(V"
P6F@)B$C\"N.A[#9AHI%%;# 0N4&0%PCY^D414J^^A'^NYD,9LDFXCVLYJ&Y@ M^1
P$07_,"^@T?[YK*?2*ZR;$'6:R0T)5- AC,Y@6[D-:$B6D@@[<V$FB=$9-QDF!9VI
P"&RO+"WD:,!SS[*Y%T3J#6;'=#E;Y 7/&HFAR6IY3DPQ:U*A!<X)8.8!P*ZW #O,
P<^-V+%UHB%@@',, D2PA"S%/L&:N0VU!#H1I$;[R4#\>:"ORQ3!X+H@*[U=>::-1
PS.]?M"M27G.:;CEZY&8:4>1/Q]EE.&?4#F\=ZF&I!6MP>#4'N+$8^137>]*T ZF?
PJFVCQ4#_SPA\EB*S#)T+MYDN59#*PRFHZS&+,@UAOJ;RE:>4]?SRG$W+U/%S?KE2
P^;U]L2_]8WQ%"TY?T'Y#M_51(1NU2<_Y6'5G>&$]WL(0A#M009KC!?1-D17B(WTD
PRRS8XV1T6\OF_/+4A(,.$)H,=K"]KBBQWM'S!I6$6Q00#R:%,[7:"4ND#[P=@=^!
PU_;4 C*:)*HOEH]\(F%<=4X\3Z3.0*UDC&@2LD.,;.=0(J0^O^U#QC"=D3#!#1>+
P8X7Q:KANBTAM>Y67<S1N/82=MP>+?ZEEQWG!M_\K14.*&?*$U(=D99O<!VAKL.VZ
PP)A-0-:7P-W"&3@O7W@ _C/+V\ITZHLN$ I]R+2Z?E2HO,U$J2*<0<<628$BL:_7
P<=4S4$TZATG,7*:(&)=@/5&4FL%?ZFJ7-& NX9R6N75&1T>+;*BH;#0;[D^J9<?#
PV^.9?HNC2I#"8K?,#..81!XC;[6CD\<N1?ZC/K>QJFF9\<Q5S7:">M8$RI9SG)@*
P1T3VY)AF &4Q?X3WZ0JJ&;E]6NH0V .= HU\\IZU2N[!>U)9V*<Z+CQPJR14P]]^
P/Q #SV+>ZQ_ O2:04'&DAP>DF R2;8,>YJ9BOQYQ$=GX-W2B?>JG-,5*!OM=,M;C
PN5KM<_ONL[7ZMMK1,H<0'6_T67894-O]UHT^EA@+JOT)(HCECXUG:B,ZQ-VF+F3K
P$7D].I!J_ T4=,6-JU"0?)#:$2*=M40_6F4KH314TF 5]O<1?.:VF0+Z"CF!'H3Q
PIHSD845!?+P5P4@S%=%S+:\&  L*DK*54&A_?D9 0T:  ALRVLMDF-$2$SP(6]&I
PML*VKMUBI? U(7F*>8MJ=^93G%S@$)]C)2]/I*WI7I<\,%CC'4*\7UR,$0<D<PXM
PKY?P!>R:^-CQHI'6MGF   &/\RBM3$[A:\SXLTI#W,]@'C(>6N.#W;<>8!#X0P\J
P!*\]).:XLJ$5C[F5RR/&L)K%E"ZF9YUJCWH:'\ ?(K/OZC#)=)_-&C//!JDZ:^=N
PP;O,N4-<)$.F5Z]SS$*;6)J#3]@F.XY1ZN".0L8R-(_6J@KXC^IES*],.F.V<O'P
PW\_1=,Z3V3>=MQ;TLL)#[ 0X .$',@+0SI6(S=Z,.U;1+WQ:BY,P>)):HQPZ5[=5
P-WG'.Q/G X>0F"WA1\M/LF]H"_**<5(SEH1RD+<U>#HIB[<0WCE$(#FUU$T[ZJ%*
PA9D=8IST^;[(E;J2),MT1]@2KBAV(F!(&:7W,;,RO =_!\4,E'"2_Q@FTXXL$K4M
P^2J!6"/G^L2$I)ZB+!C^&%;@NZQ]HUH;[B([%>\2I,?K\7<,94H/^H?BNS,8[W;L
PU1$6>!=9B((NM!;&K=BAJ75Y.]EZ3H%L>P[L<B:I"16:UU[@VT>'#:QP) 0J>+(Z
PO\8%#@)J>.1P12 .2( !ZG0+>7(R?$_[&2=0I5KQS4H&-'-@/_;[GPH%(NK,KSU%
P:RYOJD9%^>Y5_6;D^4 ['KW OU[,X%*,PZUM-5$;VILOXD-%N .V6!V_7,"W=Y/#
P-7\8SY"PR)5M'#/-R&5ILPZHYM98:DO#7L*]W<7-<_<;?I=(G!VQ_NJ!8L]$V00;
P17%&LD;"<)@"!!',*,'LEUE*[%!)?Q_GCD#;14,22C-B<TA];2[4V3HV.@+KM'2S
P7%.ZR=A!+A8W>5BHBP*[9N?HH8B:*!Q@G).\4X:/R7O#B^BWL+NP.KH.YD\/RW_:
PNI?<^&5^H]91+T?-H5V5#B$U4]?@/99#4EF4%QA44=KWGL ^$9H-&&]6C?3UE!B"
PH^O>0N]+-"P6TW$X.'_P7WH1E'502A=^5W,UX@#ZE!*V%'T1)P [_[C1/1 9DCY 
P57 FI=TY=Y9I<,<6<+4%AR6>F8R-!G93K(D*([+E#S/W]WU!F-$VVPM(J%=6%K9*
PL-]\#\I2_4G:;\Y<L'>']6_8<R'>-[!?AX YQDDD%#0L K2ZMOH,1X%:V*P<#%;W
P1R91G-91ZN2;V9D7!E-+Y,3N75"QS/7,>J7:KHMV":E E*Y1\"<@+)FL%/@WS^<*
PZ<VMQX]L2$?V'+@_NZ$T%$_#7:R6M;F5J/H,F+?1<@X-)*9[L@([LR8";8!O>==Q
P^TM ! $-![%\T07S!5A12929V'  KJ,6(FL3%X4[=@.Y(DI-WE6Y26JD7F%#2'S1
P][^[TO3I+73,IBLOP#UV)G3W(N;E@L[DVZL8E[IT89"^NZ/#EQ1HF_UY>X2%S6U$
PKTZJC?\Z\!-3-K$;[DQ#A&;E:-.#]P]NU#_C<! *[U1Q_VAEV56T2O NC;!"*#JG
PB56;TJX4\-A08$)<L3S\^<7<;[6 )9E@=AO%4[9&O<XUH%/L*!&>*P9H25Y,R!LM
PF_:\W!6$!$.B#AOU80D)E>MVI(&=.^1GK[B*C!%Q_OZY+I$5A$9XN4PR6T5T*\D1
PC#R"]!:X(JM-CY,;Y7YH4P+35,%1U3EM\^M<TDQS3""^,DT:I$951N*>S=LEN89:
P(40W.ED&<I$4BYW A[SO6P?EV#_B$$^\2 ?P,$N D[G'P4YNH(;XHB>F7T#-U/%\
P6GZ#8$9/]JE?<4U6!;[E'W$,>4@6Q,W-"YV!-+C!QDWJ7>:>LN7D*7**=6  7Y3'
P%;V O\GMK;4+F@51SX).!S$S5C?=SWB\@8Y;J-80!75K?#1,S$+,%3.->Q4TB8Y 
P"?0*4$*$LX2Z,7%:&+I\[?*V)^W5Y7Y1=A +9C82>;)S?R),VCRR3BPYEK"G6CKQ
P*&-CF%97Z-)AU[HG; (]IJHH-,U$O#W4P8Z;X.1#MV:<?L,/*5FBU% GD(F;333O
PM;VA]-^YS_M[T$/5&!S,Y;^]]3KWG *YTD@<WSQA<F1D0(I8U?(@0(%PGYM<^YKP
`endprotected128

