// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Guard to prevent multiple inclusions
`protected128
P_3XQ-["F[T#96HW$17 A.'&5L;IG /CU>IPL H9P"4P"9YEN]UMA5(P(8+70K@I7
P(4'S\AUB&=GRTA))U'S$_4?GR$'\;48EL AI_9$-I4KU9@@G;-,NRM-?K V9:V)R
P%"5>H?*,2)4+D2Z[L&C,CD"2(-[7&,U<$04SC.O7)9]AP9% 6J>COM1TM/YJI189
P!A ^A,,3TUNI46)7:@TCXHO;>Y[-] KZ*2EN.=1!0ABI+)='$>4$/ X(O R-;S@I
PQ \V]E_I^TS)!_STW.;I*!566?5WL-JBB_F#@V)JPNIRD3/R8$&M&EQ'E'6.D$D?
P;%UP'5'ZW\IJ" X[?ED_5!F6@I 2A$G3.ONK<^J>RU?,@O[B[&D+:X3Q0C(-/B_H
PJ2>2H<$[NZV/Z@&4$Z9!7HQ!W-&V'A8J3Y?.EEJHOG2ZJFD4E8=\(65:VM(L_1PC
P=<_%40W[*-=%Z3#%#A/8"I4AU.@!UNV_?);V7S/*V@6T@;"8,7X,>@],VU=W\&%]
P)@(JAT$+-,Z/0-H"/V1.2,HA.L$"AC0/B)WZ#HYW)V:!*&US1#AZ3\*@44J0:MFD
PO!=>$>B@"F;)HO<S@M2 05L06C:(_HR0#1U<81ATV8NBA"777+"?KW5.'52"<!R?
P*=![//[W9;H CQ5#32QVX;21&,\_RE:!0K&KCAW>'A= AH^_PLS=QZ]Q=@ZO83V>
PF&D>#HG.G:\US_"'1]U]P"'B_6(8*:VK(>(9 L '%YKAO$ZUXJM4/ _U96QBU5*1
P?#-+#<XO]X!6(8FUM%XRF#XLA*2_#0 K[P#LX!P66CRI9'I[@'7?I .42I>EA?Q-
P=3K69P":X[]@0X7,%Y1!% XM7XH'EY_!'\>\F3$]:XV8<F"#W[1G1=CSX>SYDS4L
PT]+EX#V9/LLK+K<#L;^E5\V[70YL]<-'U,Q-7VL%EO,SGE/E#S>VQD8C_EI(?LZ:
PW>,_!95[[\,.!=)(E].=X'HKR^EXF_GC5CPQ"11M$G#0 !V"_@BIR1&[[7'HJ-;U
P<DG!E'N+_3K^PJR=#>_J^!ND+M+-<,(:$-(EA8#&^<_H"YT=O*RO+J1$_7_QI_U8
P6U'7/X0@1+)8-82/AYR!)E+;40OU_?W IEO@)&Z\XS:KI!9(:Q01V&$&<980>%D9
PDU9[$CFT(CK);X21?6U@)7GR^VG=?.-ATSAIXO;";^QQQY!4)@NR2ZRFH,?9(D%%
P?ZK07+R%4F7?)$9-;2ZJDG@AWU)B9+U3PKH4G+S^+2,P36U#[SZ$TFF"]'A_(_@L
PKUJM ^'0 M] NAL%FJ#I BQWS3]D#<O_#QEP+A,SLXM,XRCVTD?\\E)Y3G9E1C<C
PQA&A(/P.D[>)D6[[46\8R;E$"1> Q$+6+P;OC3JR*T].W$FQ)LK#@7R%X)F%S &T
P&BGZ4$0-C)J4GJW$4SJR94DL:]>ES17?.5;EQUD\$P!R0GP%PJ':% I1XL_W]3@:
P'&J49;0&^^* _FY5?\8;#/6L+>SDS$:3(E!Z2&=.AB#9[1UGJO?1\]P1FQ8+,,@I
P.W-/3"H\O @<6%G?VW]0IC#^MCBGV/QA&_#54@BJJ>8Y_LDL!ZI%G(+1(]9PC\3_
PF(WH/&W/2BNDGI,-[=(K[';ED[$G'\,BKF@28WW*^@P7LQ<# N"8Q)K8@JR%CS::
P=;M1[\L_=I208Q^KC$"_8?@LO%]NKB^?8NLQYS+]&8*M^L;X8S^CEL^39.(]D#)#
P-W"'4?W20!5,XDI0T=9,<@PXCA=5I2X@]'W#L?<VF??X]VO5U(]]GX#&+JZ_.@MR
P?4QUJQG?:S3,8LFT&)\,6>T/C+"$9 \G(==?K+$;B8O/I"OD?+B56*$0N)>WZ^ V
P)N0I;92?_<$[ 3(Q'6?[NUJGL*PJ*RQ<RB5SX:'8?=P>AN;"M-BH?3*6OHM8'5'O
P[GB-N@7 E>6G-B(*K.=G-/>E+@D;] 4%<(!WJ*$>C\2VZXY--F"1,W1LT)]B=YV"
PC=;0$! %^J\,_OD6PLDB1 P#0QVV/011^R)B=SH%^YW-:Z:N;-[GROL=E'IEGD%#
PC36VZ;G7K$KCDG>X]K9 +$D,7+?0/["X\*=,V;](6U*O)^,ID1E[J'A.V-+'<<UQ
PZ]B?U^,,4"_ ^OY<<A/18RBM.'*G4J2G<P/GP]P3:I[W!,4BOG8>BHGK0=AS@^//
P;C\X)U=7,ZUF <++IP"%M$WIH@4S@5"WU8TO1<G*+ ^D7@I4(INB5&=9IX+F9]$O
P^C96DQ-+0,0E;&UH_<2NG,=;4X/Q:2/).[:AFO E8UD>#$UF2@TH));<3_DI]6Z0
P9X5DH0;J!Y@W\.^91HH/3C N\13U9->?)7 IM_R)H5[2Y;03#8QI2_L;KZ-=OE0@
PI[J39\DDL=OPQ>";P*;V4G'5(\"<:/&A"-J3($%W,$=F;$BK:(C[2WN ]]'Z:@2?
PDF"V@P(_Z!H4"Q-7%>XT<"/\X=\Y9AM_/Q(E0,9T90^][F+.>K_JP[,8?=,&B@9Z
P6[IX%U[91O?MDU[<KJN>YR2&,1P;1G[648D7^&A9IHA%*2;L_"Z%[PP4]?OPI9ZC
PE>Z!U8:F :R_>*("REC2&WV)"*-5@Y<"56$UG7YA3+Z=KIP:]U@$@:<;BCK;*DV=
P;MD$AD%PSBO\;&E0^T7$=5I YMVTBB,38\QCN-_+?!H +I6S I]8V(MP!ND\A"P'
PJ4QHB*(%ZD'XA9Y+M=G(@YX$^0=V>A&?\7:@:7RYSK$IDV\N'KW>N%!;Z,;_">?S
P4<.UJ0NC5(7W$!T$8J_"SHOZ=7;5-&NUZA$10'/ F*PPER_C^T.KW 6MF,('U?E[
P_OH_O1'/3N/P1_A?Q9<<.>8:5&IKT\VI>6H8NC!E.!LZQ=28:5HJ)5QG*!\8*!95
PQRZ^8-);C=I(!@:G:C"FII7>RB'WP$:?P0P:2J>70&$X-236OK(;CX?A- P:;9S5
P0 : ZEUY!_IPKH@0>&K! /5^5""^16?OCH5=H'>1#<JU7VN_((LQUYE],1S'%4 9
P;L4D^^Z6!]1"_%HO<"/*JD[+E9]_C;B"+H_F9<<YW"=>A;K=%'4TU!4D[3Q)!CV%
P2D]AS\P_0($E(L]O8AQ=TO?>U&KVFQ_& $WTN# T<W%\0=-RA8*E\#=64T^CYZ*0
P@CX.N%M_E;5@E#:422K6XAD=D0LR;)Q\8&BT-\\$&&%X@;S5-C^900FHHS%'2K-8
P:"#-@?11,"%70C^I,ET<ZQ'M8![E?,I3BGWW2]9)1ZMJE]@-4$CO]0P]*4SE6;EX
PLN*?A2)TB3%L4].6,^E%I:[Z%ORQ_?ZP<)/)D*@.O^V80\OTI$661[W<X8@8AB7 
P+#F#,WEW4HJ^#S:&!IM6J6H2D^?H%6+%(T'\0?/:D4*3Y;HFL3/O.E!MC8INC&P@
P:><!)/G-8"I1"H\Y*JQ\DRUGYV8TA_!I3JXA'4F_FA8J>9?FKV\PB=]@GW:!1(LF
PTV/#)#^/N<3':$HR=)UKRG"(S I6>8IDC\::KW0SH_$Y"6O'OT%94AR]#SJ^5M??
P%/%,#A=JL'-!-)J,L:!$U*;,E&RSG*JD1AS_;,Y2++RBAVBPIC500Y(M*Y[UF9GW
PE;+\KW,@B$$H:++A&74[)I4I/.,Y@GX&TJS/[^@_%BGAO(Q<FIB&$.*!$!JR1X:5
PT\2)RX=N5M7A3_N*]6X+ Q67EJ49OA2P5-U=PY(9=]4Y4,N-Q11Q3EPK909BPOC'
PP^5']2L;N1R:PKB,T86*,L RE?O48>_@UMY^!&49FU9?S[MTAQ=DIWU36,C/8LK.
P">J"@]RD#T!XY%K1=PD*_:-,@<2F6VDJ2%F.;!UIIBA1L072<SAJ=-"@K)<GZR0)
PX$0 "@\JP^%M2BIB]W5EWZT)"M@?Z[@/SEIB?0E3W4 DE#W+D3K2M'F]B3%2^KMN
PF0E B!R$SS=-YL9YW4:XXR-<N  264;&LL.Y/C8,HKA,P786@^HD6^%&:$YJ);UO
P7V& "O'\Q_C30U/T-9TY])X5;6*PUR\]O:.TDK7V0C^[D$T]@:D4K(L:F6H43095
P@%,[W__KG-JD.C=>2]&B9CNQZI!*/@(-Y5NJWZM7^H-G_L,](M<KPL4-B 15E[52
PC*$P*%',@X%(Q8W[GEZBFYCB&Q)9O! SJ+F/,>"FJ=TO .NE /\:2?GO0_H3#PA1
PJIGHPR(8)O;!_=,8*QDRP]&UO9*M:Q_S3LKN@9OKL 2E-9>A(Z%@D[XU\B'Z)T]@
P5OI(H -RS\B<;MSY%9=-6.MV1R[]8+I(/(9<UYI@IY"WO24INRD2N1IQ .!E[N,@
P9=+<QU;1J+,X6"BM<!!#J?7M.@/5YY#M^9VO6B5*)I[=SR<Z/3F1,/&B@Z(#5A+@
PN"('[=M9MAU=@X<H$4?U8HAC=>U'\M+<FGRY1_S&6U (/SB:"=Y?%]S;J7$$2'*V
PKWZW(<=_NJ]CWY<?P2BT_P\!)&'(V)A$;&=[G87EFA%EP0,_]GOH'%3/T=\"/Z=F
PCYGSP,E:_K$_T]R-"BK].U[0V1]BG.O'.;\SQ&^7.^H[>I*JX#1VDL[5BCNAT"]Z
PWP[F[3LH_\?7,"YR#Y1\I4!=LG+F>M^)S !\+!-+X&+J1^ZO56?4I?@*O[]&%V*!
PVWT@-8S*J/MW;IP7EU NHU"N6M%S0W3!A,@KW=F:.@=CJN8I5P,@9*(/PJ4F@B?H
P=98 Z,A/G=8G+0?GN@H6QG:3Q>8#O_OO,,RCP:(^:W&4MW>"P!<O/'RR.>-,/?8B
P[C7_Y*\M3'C7:,GM4IW7C];<5M58UP8:-DONSMOA'V)K0F,C-F_3;*3<3Q"1HG)B
P,CX?4XM CD R:/C*,<8[AL;[K1U6", \'1?S>E?,T$D]:3Q&G\#Z#YBVQR>4.ML!
PK%-E%%.3,;&I,-Q*\HNGCFYVN-&SP9C]]@0/8)/D>Q!Y^_'GN@RX,71T?W_HGE.<
P"%P*0BXIAL/W7)\#CS09R]"JD;9@1D N2V26P^9OX=.L(U, /TT:G^C#R:-'8JTT
P/G/S<+HI1P;3B8S*:ZF&?M_9XH_&MAN<=F>Y,T56@:Y!+6:.A?(;.?3?4> %XCB@
PCWY<](@ ZVB=7(2Z7GWQ(33&@:G>KZ+C[)U;)Y/S\:#/)8]2373&PA33 R3HKEKZ
P,K8VLX!NVWFW&_;K-X  9.DPH,REDF>.?@W42$!/L*PMGU'=G<8MK<.CL.).T (?
PP#9;=@W/M=!%268\!*DY87SE%_-]A?9_OQ]JS-TT>]0Q<"NBP]*,T\1&)\ZR[8>*
P3[PW2>8C@M8EP?();HT'GV!$G]I'/JT)4& LE:%2._U2JWA'0F:?H4MBVJS^BF0*
P8Q<WZ9M5UNGK/,;C4%L\_/=+_H!E,V7;\(T1VA^:$S/[1TD<@5,^."#X26Z*9X=$
P^#*A[HH.Z9K1\(RK/F"Q5DP*";H:34H:N&1($\7@M^.V^=7#GVL#+@=B13(?TMZ*
P3],?[!._X/0>4I38V?)R78=;AQ. UV;NE B68I0E_R@#A.LNP=;YPNJ8$UYR63P+
P3-Q!1D(VG'F4ZPIY/QKFI*HTO]"2CJJ)$L$R)"<#P-YWZU0<TV%FLKAT^?UHQJWC
P[]R]-5#%^95I47BGR^7=Z@,=,F_>0W7R./:Y\XNK\HXP6&:J#\A5R&TJ;9]WKYY4
P_^?MOIHM1\4HWKTC6IQ;4/5EN.A;'O91.:?RT88T)-HP.8"-EYVO1L(%2Y,%_=J^
P>Q!&[GQF8\7[ ?P=E1CPZ\'H+/OEM5L%GNP/7K+A\F?@P0GX"?<=-]]Q9IA6U[6F
P!"BV/SU,0KJ(IJ>#HI'<O9<8ZLAV[4 <B?V47Q6:X8=GSIDUN<VJ K3[59)$^24Y
P^0=B9R15NBLQJ[&8F2:9(SOHZ0#JGM+G7)(^/T[YEC>,>,)JK;U*3A&ILAC#&2QH
PEA[XH1>A L:TFA397Z6PUBW9"JE)/]>.-ZID%"B+,47A(7ALB ],O!#W1B#&<+\Z
P>@O3!6%V3]B]FD,._IR,CGY4^M3R36C<FG3GSO^\C:7^:\9N<?:\H.9J4])*G-9+
PO^=*J#?2%'FS'#+*B5DW=G)W'8-B>@-F;\,);:C!K.2/2KTW"5"SWSQY1Q*@M6;+
P(KUC6_W"IKIVQ-W*>&7HW+ W5VR;Q<M?^UG:#0A]S=E ]=]>843M@U#EHJ @@A7]
P;]*T!-T!<W3<C6L8ZCYOBS?X5PVW0\GGYK?["2@6C8.3:;0&G0@^B0U[A#)[N1B'
PB/PAF.OBB/BHGD391EO+!:71+,!^N!*F+W>->'%L96LNL-P\-!,X=\6KPRU5(:S#
P)H9/LW&J7(715V.6[A6K[0?FU1Y1PH2\?,F#R42==9N9"7^_P%BH5\F\^-;2U];]
PNC(/TU"CH.P#OQK<5S7C&JC#WC49^0,6ZB;:Z<%#6$M;14,^6%\'<MGE#A<1815N
P71PMN&@@"*FL8T-YYS9GF/1 ]Y?.1"8-"P6/0P=*R;T([<1Z!^4CY\TG<?[T-2"U
PL7T+^K#,TS2 KR$BSW'S=8,=&T3FPLAZM-G?\XS4&]#W[<UL(CA##)_&"LG#@'3A
PP@?#&-)=-7!"'$2&%4"-$157X/J=@Z$)B071H=0O0M'W^@"V!.#-R%H/E!\-6%O4
PV)D2U1<(S6JO]6TE)2Z]6=4C<4PVOI^7%O=BB-<-B;)J#,A8,_C%X^42A!\$K8;5
PF&*6A][=)I/WL0P=M !F"R@SX2[R)H 9\;"E6BP5SR?$'0)D5A4FA2*Z'CF5RV#Z
PL6Y5"8RIYLX@SR6=5WG>GNGA-N:'AHGTV2?0234&Z&'X:.Q3P)2VB@'D\K*"EM!G
P68R<2H2N(/C;*O@Z6N8%=9-W"V),;=W. #E"Q<TJ9$J,_$2GQ!$/8PO9)[SQP_-T
PIQ<3DH+D!0Q B9T6*(F5Z,.W"NB_1'[-XK2R>K "?10@#HV"(S8#3%[FE;2&%T>G
PH$&OZ8YX&\@B;43N@*$M]62M!KC<L93>#5X$,14S_!E36>*DY6'E9I;K#R8:[WJP
P@#+MA]F93OKVQ6!UBF/MFRG7A<=B8A]7A7,UR^55/XGM+P1:NF4'E@IR0:Y'G\\V
P,#+[1#%&(SA")3J;_=T/0]FZ0- A>$6#'76HR1&V2#@T%NONSE 9;S['O%3+_U:S
P52-=A,=5*52E@K[;ZZ*&7/>43O/\R&<L)P.H*UUL$0)[[YA;SH*&\G]2'O.V>=^!
P<#J,I+U[*]&;IEGB=;WF*28B>U*FI<-B0K:!.8S[[)C90 EZI6BWG]=4#=MQ@KN>
PI69M,36TIK?H<D.Y1#1?S3GUK[\(877H;7L+^"=3-:P0\6"K5-1&@-$G:J1?+1$I
PUU]0R$@;.K9>N?CP_R(-("\]YG"XTJQ=>,.S2F2<$0&IBD;X>21V8=%KYUU0=VB;
P@9;,!FT3BR7U9L.EJ ]^^19&4&9SN/9NR#K^;CW8=YVGS9:Z?":"7W]=M!157J5I
P&%_F</_N+,>\@-E!P,O]]\,GZM2+JAZNC=M.43D&9[MH#T)$>4I?[:!]$9Y31^'Y
P;J4N@'.U$)/7TIO C0O$/%MVIXP\D0)8++-HQ6G^-_2AT_R.&Y!=J1'YH:!_8197
P6;4#:&YWY$A!:O( ,"TAH%/?!J4.?<YFN )D"P& Q;0QI*);I8MUO>N0FEC8W>\7
PH.-*SZ2(-->&(9,WSQ(8!3YG3ZS!="/NJAMMNW&Y0BUSA*RVV5'RXTVHE0/Y8BQ0
P0,A"!BS$!+(%7.^-:WK21D*(G'F:XV@ 3.<$.]&/-6BB%R3J,XJ*3G#QQJ=M'Q"A
P83\61.YX;VZIR7Q_S"*!*UF3[;>5%\MKG-#>$UX\1!X.52:\>)MRPU[V$F;SEK&X
P7KRR\@N6<C\XU38MJ_TVN874]Q6C8 E-@;WXC!H:8]$?#@9UEN"K8!_[#<C&:5E/
P3N!P1[G#C$&6:R =.N U8W0\[O1.,ZPO[/<Y*L<[]LL767J3*WH2B,5=T'/WVBA/
P4@\/R/LXHU?48^G]B@'MP<967DZN>]^WL3:$HXDE4";5NNNAZ=]7;8?W+$Y9B8VB
P=1--'N$3R?W8/M],T$W)3B.[LZ#783'D.J#.UAXB\@1(13K;PQ &NYR1:\)E+^Z6
PKY^V6P,O"^B*9T[G8'Z%FJ_R&?J96&WZ1'B0!<<PRISY#2SK 2J\QXU177@4BP)"
P)Z@Q5FE:<ZIFQCJWD*F;2P9%EKK;9/#%5^_5,,;G2F\D&-+<H(7&AZ7'1ONIU7X@
P-'6D<KOMQNX^+WSR%T9-7E9 XXN<K-C>;0((WWCZK5 >+M$9-J33*W<_5%JI-,)*
P-=:O>9TYT&XY'>8FF6/T/HT2Z/(NM:F_LID9XN$J ;6!!.=&\$MAI(NGIJ26'1_Z
PJZM"H\=/+1>PY."/%FGUNS0-5<WQ+ZX/)#VJ%ZZJYV@W_0LJ+0#&+5@A_A+81CA1
P"EL.'IG&,V'\^BO8#BPBANE@VW@G 94Y_ (_CH4&:"";G5640LVQD]9VJ T"? A:
P9MW^L*R++C@;);CBLY_56Y_V2\!O4N>$A(@6LBI J-&[M?8 NZ7+' V/U@#:UA G
P2PV*.DDGKG1Z\C"B!"@UE=C*/O?*;V>@5N8;W?CRHV-%<%9*+3DAKB$1]@]W4&8&
PD[X%0H,8"=]M$?R)J-4&/_"'>=X6B%S)L@9>R>\!8&V[07<=9*P6+A_9'GEW6.AP
PUHNO4L/AM(2[5]2;9UK?I_4M75*LD4>5A:B_[3\TM+4'/)@"%)2^#'"UA6H[&$K]
P;$/E'CT+<X7%5+I-P21>%.'ABB>6N6!I( )=V"@2"K"3;,P M0'(6V09R=Z*" H$
PH Y6'R T0^QG.O614WXHB=+?ATZ0I%"WZ_2.NH[<\RA-Q4)#;),(P6.GBH,Z*/7>
P8*DSN(#[""=,3_>E?X-;L\_'.TYY:5A1/'=3S,H._V@;HZK'SO<&G0JQY$(_+ HM
P.1\4_&,-[?!O:DDDS=.T<&.F"7.&GY=+31];(:V+7A;*0;01;G"0[^7%#%/.02[*
PRF]27)PAM/I62@]'_\57L1>[B9]S;$(M)/4F:^(,VQC?&=O"5LPYV7)IV-]A)XAX
P4\"O)79Z_R4-6J$?$$G_/R^G_KN).!Z![(9$>[9;K[.-\-]@*D2!GXDO3Q/:-$"U
P)CBO@?'X34X^*LD"9WD(6+/])=_A6=J17&N41,M HD!Y9Z<;@0D'P=M99FXCBF2[
P:2CY>+>7?SDZL6PR(ZS/QQ+U2IAL3VPRQGJP> N(8<2#'$C;GN"#M@26O$L9C@DC
PC]J AKC+&$^YO,_:,$MO@^D;<D(J'PH 70]\U/E]!51Y_4=1?"RP 7WX] ,E3+2,
PM!#K>/4.CB>F1.8E9W="T;CL9OD.3Q^WZT#%CW82]H8N^6NNK=(&Y777R49O^!' 
PT.'U8MSCG[%-+TBI'PEG#,#<A"( G59>]UW6NW 3;8X4=NA;?G5+=X66?Q@'K;-C
PPJJ\YU(L'I:4%L90KS*2S;3G$39G-7B')+/'&L]$@RK9,,_%BU$V\%REVC&6KI?Y
PY$M![,]BQ)O,OM5]$=AKT@;;VV>(]=]@7R-'D,?:+^"U/(/ _;9D \4DI\.%P&+H
PIA/ABE15.(HA5(G+KVA_9Q D*'B2T$&'"T^<WN\FP,L2G2:OU^?XP<X4TZYZ;')V
P\/NZ@AC[9:;)OU1SPG)X]JZ#^)[/@)C(P[_4\LMDQ>/ORMF!-X:Y*CZ-)^(N-=H%
P#S4^8>9IJNN\G#_R^-[CL"U5ONI>]H)YNT6PNS7=)<&/&F/H_32YA29[C-K+]@$P
POVJOJ!E;V!DBQ+^42 .8Y_UJ_RJO9'H[&:^G$%*J'YZ93J<0/SW!\D#MK89KW6&G
P[-KEI2W\GMEPF:U2 $Z&@:LB=A#Q.SA;Q\4DJ.M4$,J@%_?0*J&/VA@!4M8_232F
PZ'F?F[S-K!8$V6+;05F4XMTRB/9IZ'TAE"LJ^R/=AZ/7C9SB+M'F889],0]O@/P0
PV^+*CS4=U70$:S?>ER:HB&@!9=HC0J*7$\J+HWV?:)S$H" $W8;^]4TRZQ4 K\F%
P0"XC@OB]E;G08O <F*1<6D(JT/+%T-IX<S;:1H&Z[C:03L>8I0Z1+RT)6,T28HF>
P^!;\%OBS_75^W)=_YGK](Y";STTYM<XN]4<NR0O8<F)5[3(&3,?O=!R9'^$% V5"
PALO'=I4TSOYWFI 8[:O!5SCOEXI("*[;?@[Q3\V7MM5/:8EXIY<GGO:+]TVI(8W2
P$(!3NWUEYOSTSMC V!NF;9*84U<:+('P6%QA\"9G$!+PX0&7055OBEON[V\SMY9I
P5U7E&U]*168V4PF#]"ET\G"AJ48/>Z_[4,74"F67_F@V!.C\RO7C+6>-=DH3BU"5
PTU6XQRF^L;?Y$T:<UF!BQ6J:OO"L"@/I%26/46.<EY?2P1L:P]8&9XR(KGL>Q/\4
P(@V;%@ZC%"-V>>F**AT@<YOADIAI_(K<L$VE.11RRFT*K#FH$P[QO%PTO,>&IOG\
PW$,E!$8Q1[,-#&+GO;J.2K;)-P&I5=T0CEOXT"B\\OR+>?P9$C/3AXWS1IEGDQ[9
P2[0!EN 1II_[*[MI8[F&DF# TGX*,798SJ-31Q0?XC#;&N4>@<G8=F-D/'2@?D:F
P#OV0Y]]OHMGCN19H@;,+B'M<'YXQO"(S-Y*V.E%N@&PXN9[KF)-N&QSR26U)ZD,>
P6V*K7! MGE.)H/0PY]WO0X.P(OZ>*/AP:@^=8+!2C][QA3MKSU*L)5,&DL))X+3W
PA_;8"0Z/MR=&)2?MRF3U"_!0S!TGN" '>7O8&;LJ""P"88+=K4.)+53RMT$SJP0 
P6 II#K\K<PR;5V_P8^CB'\R0YZ5 *5=']G[="$/WE+^\51N38WA1Z ^#K*;?3EU6
PZ_,Z#X^&Q!&9@6P?59)4+@^'/N5RO6]VX'0ZOM"-[QJHB[4I'?^7W!/5$.=6>'3:
P0%IPJ-+/D:J)>,9;IQT+X2/<MY3CPZ,JKFOQLJ,Y*_?3\7/4?!C*GW).4 <-"7DF
P.$!9'(GU>SONR(;IZ?:Q2W',SSQ$7%(@A6B*NY QGG[Q@$UVGR#=7F.3-N;9+SJT
P0]S#.3V68HDZW&ITYU(N<,:[DR@.IS&OXL"* S.IF8B3F$' OL77^K?/'2('(*68
P@4$@=S%,4K,2D)C'\5)M)*M\3\<I%P)'O3$-/'\J!9)"8.9BEF]OU&Y>D2.([EP1
PL'XP\<R/@I#(V5%=<"7GE&:$P5*UD?,:LWO%)D%6+'SDEMY]GM$PU3SQSUPPR&6.
P:E5UAI5]E9V3%WV<94X7H/BDX#ZV\WT/2^(OU!#I*IC,S6U&4'C_O09J>A1_JTO/
P;N[4:<6+B!M],=TC.:P?#Y&T+EOJ33J]OPCF<JV/SOY$?2U.SQH3BE7*DR0.&!YS
P8)%5U(\=R_(@ESUB7M.@N+7/==]&M3BSC!4&'.4G?(<<(TD/-X\Q D$/<MDT.>/W
P7B":U6N>QD6 1P'6QKQB77^/D$"2HK[<S'J9%,/E<ZB"=>M2H>O0[=:66X=*2>T-
PL,^-0I9N9RH-\#AV66DM*,#2FS!L;^J0659A(SSBO3YZ.+J,L9M%M=\WU!9FZ"6Y
PV/JO?\!=*!>Y/"[ J9@(2QMJ>L^S12!%A:+@92!]ELV? M"8DZ,/6)G. ,/=*JKN
P$Y*W\)\H7?I!B<5<?>]^X">N?SO$H"O_'_A<=N1]3OW9W=6'0QXYXN[KD\"CAO62
P)+:R;/%5<'!'S.M.#5;I^:OG>7!2 [?)C1MW> !F=+/-%@TR\%-92O8PFI1F]*CB
PV>MO5FNT*\=FN<Z-AY\^X_^-);@W:V.+Q)]X9X3]I.D0HKP\10:;5 /2&G/3UF>J
P\HIB\^Q(2U2#EL.D@O"Y6<J;:"?>I_PL*3[-7B)X]S- *T3R:1X@-S"-FMY5+-19
P^T!'<VZ=@_/,/2K+;-9O\Z7_(!BSS)<N2D;@M 5KG<CK 4U W/06J;(V]F>DO&:6
P^'2Z-M% $<0G+-+9E7G&_<#I%:M#/4CYIH @3N.!Q#!W!"%[1C7FTHU2CR<D9@;?
P%,PZ+,P?HJ%PR:T*=B P$H=@:B.9\%5&A>Y:?O.+GO$L&;<F+L2$('!XOCV@ $T9
PS+[#1;HZ8=U5@A.!$KI0B_@--M1>U3#]2@5-J&1@:!P3$G\"EA]0/36MD#=N'H;Q
P0_]'<AN^V,,OFNS (\23][DX?FJ;[WK&[$ZX:O#AQOL^*;BGX;X;$FE^M/1.PGE!
P/<,9T8S+0O'Y*DUO-QC5ICU6!E/?+<QJ2" V17$ST8]BK\I8VJLO2")O;\*A<>_G
P4:--=A;WT)>\;*(,5LJH4]ZH6@.L-%>.@D[D]9G@RJ)"2-!@&H7/0U^%U^*IH=D%
P[]0-N2/1&]O1[B8:N.U;B-Y7!J*7CR1[3+ ?2#7+'^4VRH4XG/D&M"LA<YH"V8<+
PA61>O.RH)*LNB7&:V%E_[$4587CCJ9V^@<K'N@ YJR^]Y_9H(V&BAR%#W;@^%Q4$
P18CGE!CTFTUD6K 6J$U(TUB+9_@!'.J+VWRR)T];H2<NHWCP'A E<^N^.93,6H-W
P=(CAIP%Y?<-VC0K\*175P6!]^&/J1LUR'8.SY"6[D%CXSR-/;T_' ?*6KG%BC.VJ
PDR@C"8C_O3:Z$13]1='A.1#D:I[E4N,%CH5KXA^4C4"T3I<'!9-1QDUS]]DOR!GR
P[T$';M0QD!C5E/Y@K]?0M8$ :BF/Y0]NYTK91MKA(Z^ZVKP\8SIVFHT_A6L($2HA
P!Q"I3R4<IE3*#7$Q?56GU)<+JO*YMW3:YYJW-B;K0@NP"*O@])TV,Q"K?0IS9\&\
P@]'<DU7PP[%5=1P7#,"#OSE%P\6X9R7V$+7IW 1&(L=-6X6;AZ41,6SRDOL>UK_:
P55E"*(H @5P80:#'\841J<W4B=%D_WIPZO?.\U2VJJ_ &,2@%X*@2Y"FJV!O-\PC
PL:7BE>17>;R\FN[S:*5S_?T:5060/\"[!"X@LE;G@A2>!&Q20Q@J]M13+8WY1'K9
P+X_GDO^F+V_K6E)DW^+6<7>VX2F99A,<\'>",9R-&.(08D>*DA</YA>KH+5$B8J4
P]A"[**HEQ:VD>#O"I@  %3KKSXGK%&; P!_OCGJS'EL-WQ^2TI'F>%)+CPJ!Y%YN
PB.>?=!_IF;X.F(&W'Y^F7UT1*LW)*H4O1G#S>+ZBAI;]1S:2ES'OPM;7*1-G'NIB
P06F^WWI,BXH^%6FJ10G-JYG=U8[^7@C'"=+M?&*4MTM_&:JD31@5D1#<JC#->LB+
P+3-7F#E,PZ%-/CH,,:O+U L 2)\);$]@OHEVIHX@]5-B>MS#I-:9=;I6.Z4_,C$V
P'3ZJT+[L ZAY\!L LH'94K('#RO@SLMO,S&D'_LJ4KT-9ILY.RR<,=K%$.HOE"+D
P^\U\G*L.($::!OTE5A?47Q=V%;D4D'HHQ6 9',/YX%! YRM$#^#*UQ)2EI:[\9+>
P%1T?%=!WT(]AH:Z1TD%^78/A2</P.ZM-7>VL$L5[%YT!P3S6L!%QO\>%VCJ^[N(3
P#<;QUOXS<Y]I)*W5*>L59ESEZ2.=?2HD++&H*]56IL6?OPO]/A!#2AWN"FZ^PG'X
P;1Y99*4&"DU!TP9$AOS8:QI.F+*B>-3F@N-V"4Y&Z'\WBQ)GS:E\U1D/Y7!J/E;O
P=2E%J'[J38_"1R9V3C_,(9!>1(!?.99:3  8:^I'>XTI^N*;G+K_(F:NZ8JARC N
P5U8IC/P8,!]>AVR]K\$R]JA)N(<OS7P["DQ%R.)Y!6[N(%G'7OV(96B:K6L<AHG/
POMZ(XAUX =H\T6"";81<6#LQRC+@E"6UGDQ#EM#GHD8K%3COL4Q?CS"EQ(>OQY:Y
P7L30T-M:]SU%03*,1G+2Y[H1\HI..25R<J#/Z/F%U=U:K71F03VQ-VI."(;*..(E
P'%)U]GR.$;HY$N5NGY)3LG[)+]DYWMRS*-G4F]K,@G$.!1^@0F!*K%?Y:=ZU07=&
P%D( *3)J7 RS/ J:^_/,$G;X<AJ^,;UQP>M\L2O_.N^O'13/<2>E%#W<"5<B%<:/
PXF')0$<O@6M;)_3_0[TKL3[?!NH"Y8S*((\$AJT32Y#VRVVHBX-PYYP=?4$X?3S/
PQU?]XQ ZUL06R1P8WU3%PJ[$"#\OYBOE-[G4N\'*]I]+M;AQ 3%&C\,J(U_7^J#[
PGJ3'].8O&W5KV2E\LN28@EA\"F[<P#$PS]6IN5-F#04AA.4CP7-E3'$'J0Q&0O"W
P&4)J H]>[/GQ?B4G4Y^7\^>%*X@NSF0;)*I)C,7@(]5G'*X%Q13N,76EUUGWL,QB
P^I4:P@C@[)(_!$VZ ?JM;!&-9)UFLHO3><-%=*#GK4I$$<:#0L)QD1"/(J.^*@%^
P?[6*(HA,=*CLF/F1(B<JQ&PAZ9DY \V1P*L:[G)G?UAR<I0 /OSEO@]SV8B^CM++
P6B;&U6^N(C-^_VX(0Z27_SG@)NFL4P,7N1A.&O!?[X<[2#U)V" WB$NN_Z=4L.UU
P OP1A%E8481WM>56YGTCY/?BOI5.YI@VA;G#MJ!1.+G2#77F?O#HU.AJGP]8GW]P
PZGJI@2=EX/*$"$6FYG%41?]Z3]4N]P!C_MG 3RE8RQ,JD7N+6*PW759S0ZMJB=EF
PE\FD7QC+7<'0AFJ-^3N8+]]!B:T/-!%7Q72N%VC\_?,R6<*RIXDG;MF+5($2E^"3
P[@^MS)PA((>UCY54[H M%&2Z[M_!RQY*/:MHEXU^T5VDITJE"[S%2?VC4!40TY&+
PC9D 2.1GLPVGZJ<>8CS16W\R!+)#:^+Z!V'='Q!Q=N>47';'M]?Y#P ;>T\=?7T8
P(4:%O1-+<_RB M#W(5(R0W06-X%;BY,UY4?@O0J?];6NGM,#_JMWI&'#O%3=OUYE
P7!>F&QS HAU9HUOQC; 6''/1$IAN@S$7M(/IF<4BM-SF+@$?,7&4;#?%#Y)%B3U/
P<!9T&KLL*,]U28A[\DJUI"H"0V\(2;SN82.+C!P'#QN(MLO/\VB,(OOZ*6^&<XX?
PO E_*"V^F,&T0[ O"4P[?K]%2_-4G.W/0\0,RZ2%\-?!US'G&0^'A&_3O_>BX*(N
P[2;VQ:[/&)$P _BC5DV)A.$_@'S3=(R#J 8OG_?F!;F<H, Q(U\U9#'**D;M-L'Y
PQW7ZBR#W-<98HKJ1),#D#.:L#WI\UY[)*IV&^OQVMM&>T\= "A"1Q"$A -.;XHWI
P]MUR$?M:RR^Y$Z -_1;5RG*Y&W3B.S#LHN=3# 4S[ACQQJ\?#9OM00C!Y?*'J6RA
P?J].= EH'_4/JO\/F0#F!(#N[Y?<K2$I)FP>3Q-E(KLN0#CO.XOP-7TA@R5+2UWX
P0@J)9I=&,CFY$@$5(><<VKER'W' C'4HQ871V*FK*0H<![QHB[?EW'-/XQ$VIO&.
PZ1&HX>.D&G0;:H'10XV8-RK%OJ+'GY3X\:W7MFPRE5S[[G7;2+T/Q+;C1(&$DQ?L
PQ?.FD7Z,JM#-K\QU;E#Y(5?VM!?+\\I[1(W+.DN'# ?#OE>B2HD#')=UWP,,,W-9
P0.!Y,"&JIBX8'9G<3.[A4V[H)=K;-OC%XL V U0]N_!4O0%-RNYL"= SE<;$)++A
PQ;,K#5EV:<?F XO7(G];"".?=U.9P'OU<#^VGH3N7X,+!&,85DDX'KF;AQ+]F146
P4KZ/A:GY,\SV6@3&)I%3.:A!<,9/;!4Y;EVBU,L[CQRO\C<])EX+;28+<L3X&9<P
P#@4G9>1KE/I=RI_7:3(K@K<IA7T'KZ\\MP9>T("^](<><Z]U:RVZ/3?K7M ;33++
P]+CZ B$"\XR5'U"O_Q,-FTOC5@>0,FP191YWP;0#,L7NXE;Y2QS1LKZNX/OEP_)N
P Z1A75C^9XIXM:0"=*>?/5>W4FZZ'6Y5]3WU;M;C5VHM5C>0"/O]7[$05%#>\!"B
P8#SII<IU;A'(!]:O8#-[@Y&B1OQ$+/NG#3[ZU(.>^X(]B1>,O\9=61/@91V&["NQ
P_"4+42NV?5B]-CN[ZS&2L[13N7<H1WL87<ZC45A8H:V9-EM4Y<4CDLHQXJTZQWX,
PH \64<SZ^.1!HCYA04 %=]VKL!MMO+] W&3O:%!FE2I-LSL.]@C=@JZW24OX09[R
P^-(."0@BCM>($\'F,6DW!# L4^",F%3\BHB.P]^PN3E+([UAE ;7Z:?.J.QH603P
PUWM;YL]^C)"VUXN*K&0L !+>MY_CF.OD"#A3LQC%"9OJT7&A+Z'M ) ^UI^WAJQ/
P/RE29")ZYC!F6LL#N@+PD.5?2I>,A%8( -2B^C-5X(A"/?7=&MRZKLGIQY4@XL%R
P!9Z/G!UYGZ'2?!VSEZ29.O;/8-U*D)JR.\_\=@7F3W8JZT,PV$:R6:G&B^.<]5RL
P5+%VD^\,G @VA]@YZY"HY7?Q?5L>\MM+(C*)6]X19T^NMH@;L4FB[W 5\&''#FV6
P-S9#4"X%]0H?!P/ ((4LI3)%Z'>_\X\#PM0=*WX"=I=BW</*KJG#P^$&']4T2Y<8
PLH3 O<>/XS.$73>[&^]P(DQ2CR9!C_<',[[]./4 4T$#D/0=%DO!CNZJOIY/\UVX
PGJC5ZME($+F@[^C*:%3\V\-M<N84JK;O+6 I-0BK.UB,)>A#\<E<4T#E6OF;B[6^
P4N>9UIL7L%6J]"VF>GZIHE%:6DFXHZ(M&A"@,5N8+29>=90(QP,&S^.]42\&/+_6
P:=6=3II[B6CG[/NKT;!DGFX"/D,?;R;">1'+LWOFDH!X\,'\\$1@X^ QV'@B6!'X
P+,; [=SN1)Y;"H):5C8NP%$Y+DW#+L<#V))P-PR%/&UDU,PCQ6NB_;,\%IA0JCZ#
P=O=.R\O)R$VK/]P&%(3FK0T2",Y.M,O%K@W3 F((NI(J3AB@"7XZX9%/P(6X?<O"
P#(E"-R'SJV.IZBO 4Y@YZ)DI:2$D5Q0HTLK$>+ 3>*:B7Y8TVQJHLP9<TAQ91MW9
PWU+![DR\\]J%KW&>D&[ZZ+T&9&1PPX%C]8:'KJ1*EY>(R/P6C+4?/9N%O'(R[L!*
P/NZ#H#U[%^]2\_IYYK,U8X&-SB,S<3G=5-V9A6A8%F1F%38+(G..N*/QEE*G8B^8
P@!)]J IO5J@] U5S=B:85H6=YXI+C;O.%5ZT IZ@(OZH-[OJ/'?&PAGFJ<PZEE68
PED<K3P,)&'=*3VZV;%1U8'G=&K^PF#2MR-41=UQY54%IPOX&@O<%%HJEWO)KSK]L
P%00HAB9T5YG.J-+4DT1>"6&M]1<6XR7VZ^-;8_4-OXA3 R+U<,A>0AN]/<EBE"R-
PM4TZ 1G(6HGPXZL/PZRV$*O",?4+10A(58V*%**PJ8&,M:E9AR)*[MAZTHBKSKCL
P0VV\")JZ+#:(3(I%;+-0K1C2-M::( #]\^OKTNB'*7:X=ZZ']BKZ5K]^,T]LVXS0
P)V@8^M#]7KHST4OY%LQ9&3DIJT*4B+"=:6?R=-Q.UG%O0O@+A#7UJY_8?OI !-A&
PX#=[( GVM%(K//$=9-R;1>ARZT[Q^3B>S>K@H*^R#-E.+!.ZZ;=H UHS&6]]<=P2
PD56L!Z[YKN@6& ;*[)-15"I+XZ)JJ'F+=(;?69VD<E,O$IDWJ#O37HHDGQ7G1>XW
P26&%L"S/K8)2&7A8 ],*D(B2H5-/<&8$B_?A,=P"EWUK]DJ;+O^UE-O H.0/_?BO
P]V47,%&#">[.4\<'7!B@&>5  \0U1%V>6SLE%7.M!KU8WU];)-@/"]2U_Y^@Q>><
P3+4EJ[NM5_FU.CTGIV0\F ^!WJI/I 89K;U/HGI.2/0PUZ"!CJUSH-F[5@,JKBA?
P5U+$Z^LY#SJRX(50[" NH<>U)NGI%/P'DMR\P$[>\<DX(6P*>UZXUVFQ_J/4BIX9
P\++U4)@NZ2-C-TT'Q\38.TP0WXIY@*/RAK 72(?*T40PH%*.N-7!'64@$F4J)JY2
PQE=]Z2]*O: #T?Z>T,<^LP^*_H:""?U6*)0QXSV;H_H'X]/,BT&N8ZZG>E+_&)6@
P M4-$*+DV0(-.W?)C4#UB$S?(%WZ*;5\^_V>KC:%$(P;>Q6#,SW5Y FZ%PSNY_.I
PR*P-7%U& &BQ_<)>W!IX(\M3N^SOAUW7M/O*#9)/":+G-JLM1F$RM117G0 W5'[J
P=G7Q6'<X*9H/<#'Z# (0[D-9FDHO!F;*7K\9O5 ELDGXT3C%.ICKW\G\XUKD?V<W
P>^1Z)!3@B=S>L2Y\F@GZSVDV^M.;H=.<ZVG7N+487V3!>3//A161#ZHGT@HR#H<*
P/*=.CUBFL)$PRE?!=@K/T)!7Y;U5AE)J(T4^9RP6>!QC[[K]XH&4&NAT*R6!Q1<=
PJQSUJ(C^-Z>7FF@HI@70/GX-@'EQ :27ZUM)/>_L!K3329;I8 &0CX(#ZM6QZ8>G
POV3TY@ALQ3W#1]50XMO4;)X/J>8T]E7!-]DJ&*RD.S7J2+A/ ^_RIGB8,>4"B,J[
P/+FW^9J6B8JNUXR[EYV^&=F@.&//J;P,&;]NXS#^>"H-:S\>A+X21IEA#N#OZX2&
PJ0S]!=Y>:*[M>& .*?\/*K17J](T='XOM7,?,Q,ROU!5H12#F>U$%B>*E],1CE.1
PA7F@&KV-0'(XP ?C+[6U!(B^+.C_V$AV+M5H2?X)C,>@I$XD5"C5><RFD(&"D7:<
P((:)QF5+CM5(!.:V=XE53-E,;<^<UW_'5VN[IRD"A(Q/Y&NIP*N AK_<@X+P Z@;
P'"B=X'?Z6["GA;.%OO8F!*?%P$K4T:<[3]J;T78YZ_6R)<*G+H*.5FLT0TIN>F-@
`endprotected128

