// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
P*T5^(../302@5>G!&,J?0/S/89%@<O.TO3PBH:S=*1<$H=$SYHG1R?MB7B@N@JTU
P CW$F.@ HRJ!>XV;J.O] %UB5Z'#V15@V80!?@UP*:-1$3#%\*@"2QJKYXU;8CKW
P2_!(R*L8)-,VUSM:S"NH(B)-V"4G.?'TN;SP>2Z7D>-8.I A[:@(KB(>[A.\*/7[
P2UW6BQ1=I=D-NA3$&+]'X]+CF$SW11+2CCPF(#ARFG@$;&DN)GRR>DP.AH4LN_3[
PA;9REM\EG;W]3^0I]7&DLN]4/_UGO/=(HJA#&Q5UIVE]H"'C$6KHL>H'*W0 3G\=
P5)X84L8_F$RJT.WX_E0PK"BQ["2IV:>JVC,(=ACUV]=-M0J%3(=K#&&&^!P/#-C>
PSL?C\EQ'X6>TW +)=-7"^H_R]F^Z.+F_A7'<MWFW\(6Z!@ 9 E6/ZE/Y8K(>FFRK
P\=XX9E!3GE&O5X\SY[!@:14.UN@+F[HTVA+9>D:C5[<S(L:6F2[:CG$S9+AVD(:@
P&3B.D=!SM2X_H1W8M&<N;F&!RGJ5]KH>WE2K2Z":-,%K_!@_X$'_SXG#PI5Z&O38
PACO1)=YI#B8]&PM^S0BZT%48YL'(V(COPX*_-V>(KE<ZBHO%X<BVB>5F9LB&@@ /
PE_L<-'<"N#/&YO B)FHEZ'#)PC'3 :1OSN7_U.K1<P$I-:LE]"*PLVG"+URTX_V'
PD^U:@SI:VF8IJ(-FFK[5YQ7I!R8>?4>=_/J@=6@/IEIO0B.N[H'F1_\G,(JCP?2D
P2;,1B+NND+$FHX+,+@C-.#Z0@IW$2_^2&!M#FJ-<X,R^.G.&O^GR&YB]>#"T'\5#
P<E=DEEWGH.L8.V[F-K,$9$2M>H7/.=AKMXOY[_6N1"L2;F M,^5-WU&$RX)(/D]$
P29GBY:5V_=>W\1OXT/_[XF%C:/9Q'4^^:]PUDVU[M@59$W%.J>EQ/S/:UE0B:P*Z
PT=) W!:NOVOZ_^M2FOQ4X](\6D45'?1RK.$R59W"D++DH#F5^XM;6=+F;XT=@([W
P13/%Z'CR:?>)H8OC44S/0:&C<(0G]#S/)!SO&*^!XEH<NOM7Q89"EQ&O 5?2C2 /
P#4C9BEJE23'FC[X21Z^45'C@L-R8&*Q/)1&33&.MLHV88.]9,QP-D7NW);SS28<1
PWGR5T:.?#ZE&K[JIP-0:=!6BR;C4?MJ3V8-W1S2Q4W-Y"UL])!>!R>!L"11B,\=:
PD^"A8URDD?Z?W& .WJ:9=R!4\Y[_"F=DFYS#U3/E.X']2AISR8L'!D B<9,M0"R-
PKW2@@O-$5*IL9F!'%>NV8^-PI*A?90DLP&E1JF5GQ+Y(O]4$LW6;_Y&JN,#,>,1/
P%1<BW'Q&.TRBOK4?+(R,#1P;"VWC?P4UJ9(W%I0WH(!O3_.#VI. ".NF@B7[KFK2
P&Y-""B;BRJT;*1?X9\N_:SQ3HYY.FDA^1V&BPB/A4?<4'$HM?3+ 1N+0@])R.9H6
P(91+QB)[,M-L0,LD1N27(NV0]O3E4K/FC@0EX<$#_[_& #/1H0%O/CWFFJ#*4U<'
`endprotected128

