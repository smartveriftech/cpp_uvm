// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Guard to prevent multiple inclusions
`protected128
PS.U^H7,)&* P15FO+4GMSYF([Q7(528*\N0T-7F&BIO1C:QZ_5:3^1LV5A,&BOM5
PLHH,@HL\6FAR& Q[\L939\KXV^!"K5$^YSN!A*E[DB>VML\II<4#$'H+8$BCZQDF
PRG8F@(C3/I'9WKO_$6;A;$>5=WFS!D.4A"4@(QA:TL#EGFAU[( U/-[D1O#]LV_T
`endprotected128
`include "uvm_macros.svh"
`protected128
PQRYZ@=CE:)!LU9BL-4,]F!P/B,'-$D_?EN7M%VX=Z+"X+A!*4(3[5=!WZL ,#U2\
P) 8O.O&[^AB.S]NT4JSL<,?B%M"_[2/<>;806=+/7X [_\FB> ?G+WMO?N&Y*/8E
`endprotected128
`include "macros/uvm_dpi_macros.svh"
`protected128
P&N3O]G84PM6*(\PTP$2$:0 BP(F#6 U2J'SX1C]"!^Q\KC6F,>S9"_\"K<K.9]FY
P+F2#9_2VY#54]0'7/=-GM&B#0QN:6<,0P$?B_H(+T*H]:YJ)8+<QTF;^Q&*LY_Z,
P6E4B<#S>,J3T99/^O/8W!H:NB\V"=T4\X'H@ES7CY0"F&;VO>[*UY^L!)H,V8DYZ
`endprotected128
`include "base/uvm_globals_dpi.svh"
`protected128
P[^]!(RL=?WB%Z+>X)J)2RWD=Y\L+&>,@7*@Q_Y*#2U%K9*MW3'63E_1_?M^A(R,0
P,0ZR%\*V2.857>;H782AIX[]#B%N@WV+L,U*Z8V: $Q,#L($5Y"$'EN%\ZW1S#99
`endprotected128
`include "base/uvm_dpi_defines.svh"
`protected128
P!YO]/M33N_^.RK;#W)K:T?UHD8,+0MV^901,Q:,&XE/P+<(XP?$CQ.M;2G6.1: 4
PF]I--7BE7"=R*YCVJL*S/7AMMW:'32:ON=S:_0JYL<APF>;$0OF/4B8-\2MPK+'I
`endprotected128
`include "base/uvm_dpi_sync.svh"
`protected128
P5\A%BP=]A8PJ>S#YS0'SI,/13/V6<HZ&L]II?NQOL.4HYF$!2"6=N=_48;NO<NE_
PB1IAO5'!O<E73]*8AN!),J!L\2-[#E[YU6\-1T-@5:Y*J&<Q#;((P6<Q9&SV=QU(
`endprotected128
`include "base/uvm_dpi_root.svh"
`protected128
P2:-8KQ <Y(^@N#@C:6%#9(Y]U:K9V9!D>%PGDI]#(MA%"C>A:[4O\<H\VH;:C_'6
P[5WVMMQ\1A7#CAH^+,)$.!(K)2O.:^7J>U&_5$8TX*%+GO0;LIBP1.@H?*!JN7UC
`endprotected128
`include "base/uvm_dpi_component.svh"
`protected128
P;WJ9(L=I1OH*VDN=E2<'6MRY'CZ9W2I;P665@0!Q)JN98I.-MII%VVBNJ-0(AFE1
P*L>)\D?Z*^6/-&!5CZI'FS_\AEE3BS,K7Q+[$]*-VYM DG%@G-ZC7Q/2%8\*9Y1/
`endprotected128
`include "base/uvm_dpi_helper.svh"
`protected128
PQQ\[?$M2"64-_:H4=;NT06J!ZL^D8330HU)ZV4WZ2S#4=5+J29#=U,_;8;&VBQBH
P5:0116FSEU$S#WP\A8;]2C.^((21<Z@B+,&B(.SXTHIJ=)/%#ZNE0\DG$BECR*=Z
`endprotected128
`include "base/uvm_dpi_object.svh"
`protected128
PK0BX:=WR2HH(,!+J3@LB2Q]*CTCEL*Y%ZN^3LT1FZ N.1ZXE.BM J!Q2+ >X'.Q3
P:'-4:[HB\F:*J'*$:NV#,\ 4OI%VGJRGJ\2@XS2N9+^0)WM;)1E;-R%?TM:B058I
`endprotected128
`include "base/uvm_dpi_seq_item.svh"
`protected128
P'Y%(7?4AZ* [?WA"V""1@TQ@*?R9=^!M]C6I=RP)%'O7UL@-S#,73V05K$=#POIG
P%\B3_A^NS@S/[22&V]A@Z!A[1GM/9.>FF%=GJWS N%;SGJVF)WW)0GI_)<I<1661
PC!!D=RX';*9?51*>8_Z@F\M$5_#L>$@(\=3O5R$#""K_30,:,FR<%HVPM=9#MA[!
`endprotected128

