// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Guard to prevent multiple inclusions
`protected128
PY^U5$].]P(_?]^.>K]T, 50G%NF2DWIN*\\:TC:3Y:A^TN-*?;WY<ITXLK ?CYX3
P6HTY5XU,QISY!XK.\=*TVQXHGZX1O)$V91]AVG [;!J50"XP]K&&>V=K%C\W*9IP
P@%%,(0_^H]]^0C#OM'W->S@6 'J 0,K?-W$A,H+(&=<ORA6T]3\D""V7XB#8"!8$
P?D\4U]">\6+E>:<HK0?](4I*5"!HZ($:\IJ%,.#N/;>[9A^N<UE.T\9L)R<# (RV
P!R27@-D2B4D][!\K846*9^%H>#?[B'U[YF*7\D3:_.KUS@TJV7H@-OQ)G\(I3O*E
P W8((^?ODEZ EHT#+NB%O;'80'STMA#8%TWM;B@6DL,LG0ODJX$:EPU_5/9/O,+%
PM?HM4&6J HBQI-/]6.Z@$:K;8UMOOY$43/SEW5LXT8//HI,1<:LH1[+$DF%B-"7!
P(W1C]+D]4>KI+Y\F8V$1V(-A>,GPKV#KKBB67HV6@_-=:6"T+Q0IUQ6/7)"AR'!#
P07QQ\,_FM%@6E:"(Y[)9_8?.Q3M"SD].S9\J/80F49'(6ZOZC[=[E5EU>V[9:.HN
P71=8M;6*9S^P5]_2@(Q/?B"D-._[>9,.:8^-" ^5.E-0[/28'IF+=6NO0N(NI%[9
P3051_&"CC.8!%$;<H9Y!"+DJZT\<N).5V_X>I\Q4D<JV!^N8?!EO@EQ^1'RMB!2!
PWPWS-RT1?P8V1>6-^ E25&>RC$A80<_BA1(K*+%+-5Q=D'^:> C.T>1]5^75"TD@
P03WFK<6W6Y$98LA3;*8[H&^_&3B-P2GN(^^#-7G3LM'S1))<IW)ZKUD]]077?^S^
P<;"F43R?T,#&W=#H,QL4*\$I)4O'@\D\5(U&<IGH81U_WUBT-AR=.K]/-Q4'.ZI"
P]LH4O](+YOS,/D9A"&.(Q<M@:1]N-,4-"L6+@IC,MH.,2<WL,ONZ_<BO1!W1G/:'
PV?!([.$NIB!QMJ4!$F%6#:9A_ST(S'A@*_NI-I^GL>H2WQ9,8Y5BAPF:4,0\35E<
PQ_W7/J?<ALBF0)-I11SFT7_ ,-#Y*\-^!IC6Q4 QH>9IE49[0QEPN$LD#PSR@N 3
PI:DPM 5K8(<YC_<I3ZVVQX.O<8STJ=9!.+'B\LL]-RQU*3UVT<;_OH@<KI5Z&%X.
PR= SC:&\(&MQ[(*<7V"9XT3"N2H7&_-.RAN].4H#MH)@C1/MHP7>[2TB0*,#9>#"
PL,:(3/I;E.C2SX9:.J%Q2TU]=5ON5PKS E71_1NNE%JDWJIB'N/55[]B+.HOWZH4
PCQ/]S[.63//V2(X4T]<'5Z]WF0#Y,2;&FD?$D9 $( N<U7^MB0" @ONE%AMS8 G\
P]NOQ)I-T.U)M5+72F8U$F7YV<K8LKW5<0%2>HH\C72]@*L.EG2,5HM/"$$RHQ?"D
P0#Y4C,0"LK^G,BIG3<K\2ME,I2'->L "7\4_'I+@I@U?%F7%BW;7:EY/2J&[\!WM
P)X'(X'FRJP*A@].G2MQR*79Q^VKQ0>!&$HHJT*>L1JAP1Q6R]CB-R.[G>]<'Y59T
PF++HTAY4W-RQ061H1_O%+6WU O=WW_,F"@5P:=IWP>QHS[8?)6:TXV7&""0"S@.3
P*K'E12(7HWM8]AGY00I^*06+%-9+!94C/ZP*.>9#3UO6M7)5WL/<.A!TVI:"?Q'.
P':"WDD:;N%'^B*P#$3Q/TB3=5@7)NOL2AHF6_??*UWQ5UG0PXEA<,B+,&K&7]X-V
P<B,ZNN^V30^[@Q7MIDUUA,"G%TX7)F)95\&NLQ,Y]E/7]8#NA4<'97\EO91[-;5[
PC1W#!'; WMJ"K((0EUPVJN']4;'A9,]967:L '9)=P/A*Z@E:(!J1N6YYZ(K/9@V
P21L<"X!3(M&DYZG7EQ2Z8]"<2-2^0=7=\NFY*<KC9X1EF A8G$K:6BX9O^DH9RT1
PB+505<KM8>2O+%S8.ZI3R-%O7:&1!E;3.BFF-QD2B==WW4'#8LZ$R>2CN[ENO5*7
PG7D?]=DY GF.YBV^UH+'RS>? V!0!:@"\%K8^?C%N>3K$%R$+R)RT-B]IL_^:_VK
PE)BK\,=V -A@J%,V!7U#EDX0]RO98 $T2P*;<ZNE^5?FA=TF*WVU![X?H]G QZ^O
P]&4"QE7EW;\Q5 $VVG-:!;*P@P]T<Q?OE;4&+A^$"ZMAG(*T)<XCE% R$*)_.!J*
PC?=6!\.&UA+#]]9M^M0KO[SH+EC#T- CDBO7$FYF@@=6$(:V13W_9/-GHK-HHKJ.
P$;ZQYE7>V+X!F401\[8 '%74;JW)-8WZE?T)?B.:+;H?>\(.=E]M+Y#?RHL-Y^#"
PTKI+LC<;:IKM8DOW"&&9(-]6F\9RCJ#D05OB<L?[770:+EZZ&5Z$R<A"_DL:H:OD
P>,?S'EN$?L"8AH7;QYLMU(C%/9"ZCP4P<-#0.*DMLX/LA?A/^ZY*ATWVY& D-FOQ
P7NVK46B<!-"^D U3Z3JHDQ*-<O>:H#2O3-"_0C:^0XPWZZ8GOQ.\F6#";#V%+]3M
PBF-O@%Y,9?#6&G ;D-#G/'YT%7,\_F$:)/X8A\KCY;'=YZ&*2WHH3]*^UIA)'.\S
P+S?O*@O=4,1Q"=30)-<_%0[<U@' =MK;-1,_ZP1=^M#Z1)>\^"7K"0?BG@&I_X*@
PAC^H#B1M<3/]K9^JBLQY9J#4&T%)%YQ]1X2)K5>=\NY',"I\X;)9C!=I8,@V4=$ 
P[QG::!MYZ;4L#Z0H#Q/W;G&:F2U.[,+"%WM R5Q@B:L#<8G9UT\+_3^E,SE$<Q+N
P,W@S5KQ9A;Z>8<J?Q-A\Q)D+.UN$(2I2*+=R5UX-;WSD7!%=3$#V,U$<2K])W4^4
PS@A,+**@DKN*%3#F" 2J-+I-26$&D]IK;,A/D!](ZZ.BT+."7=U7YSS;,R5<A4Y6
P:<H&M!)ZWU%6$I 'BP*>D5\XE2GL[>M  D\$>;62XFBKTL3]JB"<YIGF,UUOYM1(
P*LRPO#V"S>.U;?\6 7"K&_@F&#B4B5)WIVK?EK7?_BTI\\J+ZCD2BIEX7W!)+UTP
P'SFWH!&+21<>@ #WONT4K!F-R9'#53#AU,* [ ?CN .1.%8W3>QV_CTVB+B!!AE[
PO^XL](XCSM6A&-N0(?9?E)W[P&UIRE[_0@#;WJ]("RG?) Z!)6NDRTT:D3ONZP%-
P6C.QN5C/,E@G4[:M'&'C8[,T,H"TD7ILW[-4CER-?L#'XKZVC50EV6S<SL,>[ BD
P%WX8_J#=BB0[8R(=NOJBU#Z_,#:4H:E>0!(/%%36Z8G4Z=A@QS-:7>5#F3S?+WV,
P)Q(FW=KQ\TE]<@[ E@#>:U?LT]3OYN3A'=PSWU;=*MF%S@8*BUJ_"]+$]M8K*A>O
PF4[3:B9WHO?\=/IB$IY7#,E>DU[+SB402KI(+30GP>6&/E'7W.#SAXB0(#9RJ[N*
P#T? #'<"_I]=XM&5& WH;9GZZDCDCP_'#/+/R'ZPH! N.R\D?T+I8<^ QRI@@A)0
P?ZY.%V2Z9[0..M)KIV7A:[_/+)OVMR5M*\GR.E?.O" N^[;6Y>SX!A6S>(W?+978
PT^".$,)/[#?LL.I?Q8CQ,TH7XKUX*.50[:Y<7/E\CVXL[,NNEVP>H!!%1>@G,]ZZ
PR[+>JR^FQ$+!EK:'[@]R2E_!F.^?B<:]V@^H:]^PZ0CD]>8MFSC[A*Z!5T39*Y7N
P@-HXH=](]W5+4:15"[/5 .G%C((5)ZR&U]!^'5'D&G*\M\C1;^=J^WNKX'U (;AF
PX;"G_8V8XS$&"]D%=Z2[]D=PS'K4P3C@X<-\E_L!D[>"S%%**]Q,J0JLZGNDJ(QJ
P)EAWO!3;]/[#$W]SJ<@RWP+CJFTN.9Y+.1&PO^_'#/1>B1.6&>!+];W&3'&F7?/:
P=7$R$\=_(4T(@JEVZDCT&[ZM_@6/Y E_>4 (4$ZIZ^,T>@$BF<ZE:8^+ (^M?TU^
PZGB=34PZT4^(^B0M1(-7X?WA>^+,GC3CVTUZX.4TFDZ/PYO'WD5JK:DW<5HU5E7%
PV!T"X5TS;KV6Z )N9U")3)W+X:ADF']UO@&1D#LT]VC),VN!;AH_4_HUIJ8D)'%K
P"=W63XP@.V,5^L!B&"[A'_U>31')@*49\'F#*CJ0I(Z4G=DYAW7979S]ME P_-'O
PDK0I<(6 ^KGQB&)[2@%S].VHFSF=]6,]8B.WF_,;.C:]^CS?JZX(QJ#7N62R,GM'
PP^BD&=/]T /[^,Q0DXK@)V54\6X?3I_=9C#> =N945\3@HDAW(B_..&Y=\)HQ\]K
P&.'K7/; HLS5%I(:/9.N\-#\FSG4X:%J8(##2UXH4EMKBY:,<$K:TZO,)-A7 ,;E
P_)<!N\Q8U%NC0MDO-2^;9Q?]PE ;($^B\>>D\;%DY3*\):#07/R+H>ZX) $T7(H%
PI1EO'F9QO96LWKH:1=Y<50BY>]:X6P?Q/!CT3'I2M 7PUBZ]S=.$?S2&] I2 SG/
P>*UU>\^;EVTMF82:@@_B[POV<EA21US[QGKX<3V5]4O;1\[,"Y]IT>< =NVW/-1\
PW(/_W7)LUAX%EZ($,*0U\'YW]!\3L5%W>SUC?YJ;MK=(&LFXK$&'UXM0\@YRM%=2
PW=/]HU.?99?Q\=M<PS+)S'=1E'[PY1H3Q(JVCPD397NP>6HZ;I6Z./,?\A^/5RS&
P:AO?283^*\&"3,Q]EZ*C0.>U_(K,0YK9'=S]8]!PQ SN4^81U<;'Z%X!69I6\PU@
PG>0) [DVPS4I7/JF'77-&.WR(5F$3<"G]D>7<R18JIL[XX3FEUX3XM *9&$8PIH=
P+U8A4/H!X"H@'-LPZ+9#XP4B( E A;K:X"63"/U7Z,R-,%!%.A=8BP11#:(XY[#G
P+):[_7S_ DB?77KC2@TGEWWEJYX\Y>1#!< \TK4Y,SC+/$M7N%"K=9M=/G2Y_FFR
PEG_$07]IS7^G0,ED]R.INMPP+]3 &'J'>%Y6'QBT;12,7_7A!$$],*(9O\5INV1U
P[V+Q4GD4E.;-4X3OZ4Z:+@^WT9^Z%G<9N$"[Q":(I4.93,&O6'%Y/*TJ \'T_<B?
PNF]KP]ZM/CN*-TGY?2XV^NBO>E_8(EY-WJD+(,Z/#NX4F?#PG,P[GPUJ7B>4$ 7-
P],;@VD'R(%[#X<)T.5#DU\CJ23O.I<B^6WLZ&R9^/NLO4?K>?C1R%@TO%+<I_]+2
P:^?U\JAW50T:B$KS=TGHZ/1Z?Z,1) )KK;?!T-IQ[>(:55$6+,P27)7-"GIHMQ'7
P/08JQ9B0J$O%=^/++N!?\RCIW3UV%DE^S=CBR?/]S=@77K:L=MTU8WYY3=:'XR=X
P12A$^\&&N<2,D #5?FYX;$- AP$#T;<#/N=L&MD=Y5'A.6A^!Z]Y_LI\6^3%%3A]
P4J4[EW@(]DH%D_=:UOT'&Y(F[4,-C'H"(<1,'TO?XL7]D?_Z7,)!A=RO9<A42R >
P9I<4XZ9D*2<PO/PP MCW8F;!?QBHU>"M<1+D@Y-]SPH:7MKZD)>EE<U]0*ZM1%&$
P:&0>NP!L;N.\L]*8J6 V!4A\/:@UYOFNO<U3ZJ@'\S!GK,#!],$,1(H&]06%YCU>
PJHDMVGR!V:;L28@%GS47*$\K/&C]<S>.AQA5=49-Z-1[6SIH![=<!4/_,ZS]9P;_
P-VIY1EIM]BLTF_ ;!WXN>R88P^E,H6O5BJR#E/W.&1:ICQ0.\JV, BXSAOXM2N?O
PE.3?[DQ3$N3&I6740'DHUHM$4.!O9@-""7'EP4T@DH3X/B/\E?:*CX[-!4XTXY=W
P_)D+/,:&EO2O;J0."@_\-'Q;#)U8]51Z-;7"C/_K*B@ ,RC3E'PO.&_ \[70KD2M
PY9O_&KS+QI:>!N7J\NR%I")(*"J<6/CTE-_JMY],+IT&U&M3KW"-H0IW3T"K/,C'
PW6HP7>^-W>);W2]DC?<1E%O_@VW/H]YEU,P4-)>PPK77<+3W]E$/5B;M2[3[?I9V
PMZU-\FZC#YX]P$I?%I3'TAH\*U%DI# UHX<- BP:7%?)")=YT2A.?\Z>UPEL2J68
PNKT>CX'S$T_,2@+ #\LZ!-;<D( ?&K\LI+Q"YI=A:?+1D@J\$:/QKQ#LI4XHFZ-<
P1!B5^4B%#8\CY%E8[\5#GPI52G-G/0URV1MXBW]4.-('6%PUV?*TWC$T9?:/@&@H
PW&%8^C8\;HQ?4$3":U\_RI)'PDG?JID1Y9"2$3)? /7Z45+,EDFMW]Y6EV=++*71
P&M,TJ(52A802X,8]76]Q =M@?UCT>IBHEYL0/?H#XBP6AR_N["OLU>%.%-F/A">B
PLGO7WQS*I+JGI1\Z<;*?HISURTFN^:OOY!6J%]H]::K4M':>RO4U\K8?-<R4$'*Z
P9@]VWO@3[0H_M;;C0!]&-(#4YF!XS#SQT WF/DMBT2-+YJFF6EMSN9]!#M]PCJ"R
PKP)K68+7(O4[S-?;'%QKX?PW%CKK^I?GT<<>J.6%S,+V'#:O"T!8[L#1LKK#@,EA
PZ=$,ZX*65-PF>R(^<98O06,!B-MM%ZLP@!#JR)U(!^7W+3X ,$(1>QGP)_-]":?_
PIN1#>/TV5=WH6 =E1(]"RWB(/ #ABC@28IVY!\Y4[1$%=JFD)4ABR]_/.2P:!0HS
PCB*Z*$58BA8<^ &8X!<_9W<TR=,//@&YH3=!&9C$F_Q%7:[Y?.Q1X/E#G\B[%LX?
PU;9V$NNI:%0) @]/Z^6N4FW]PE+CXP+DHT(M^\'F+!0<641(Z#*M'(.?_(;'83'>
PL5$+8C[Z_#1-+<#.I+TQ'VSL?6Z3E[7%%W_3Y(QKD_B^8=YKJWOW(#HQ-<$806;S
P3@T$;'3%@F]_GGX=:I=A<]U3Q'LR:%D(/-Z8648AH;1C90.\,H1Q<3K,K2 @T:V%
PX05H+?Q+]JI7P1"GW$#"6J'+F 6X"%7C!KW+5REO:(%Q856-@%6Y?>+E#G<:?,$?
P,[#$WB7YC,!JJNM51X<A/8<<MB)>.H#RD]8;O^IQEZ T[4W')SNJ*WLF(DPR;KXD
PX%$T;\3K;)KL)KG? E!^D]-6]\"%W)S7F[N>DA)EZ\8)F?QPB?+RN]%-G:P(B^\Z
PFDKWL=#,^L$918' Q.)"-\R,NT-+SNEK*M< 1P.QWHUDK[YB>]D(,P%JHDC".'6\
PWTXF7+!A,*C["))JWON")5B,R5PQHUF/6#S.4I&*5E-QVN?Y%5-^GJU\G($-Z<60
PDVI&-#-H1L/$((+1JF+MSKE'Q@3O<KL=]%1FV]._I8>0A&=77A0D\?I>4EQ)_C.A
P*I1W"7-X*7W$M"W], V/YR=)?T!HD:E[W8F,%UW\Z "9;QY\GL6O@<!O$40B))L<
PO"IXCG=2:Y@\"1+=#/%%FU#&\V[6T@ELC0O]?>$0/G$^8!:\:H7^_BAL!-,)PGF<
PKI:-/)[_/#<H<R;@8U\9<LO3XF)?NV>]5TG:*7#YA%5FJD(SC^6+=FDHL6+O2*(Y
PX%;% Z!V%O?=35F&C*6E.^NA KI*CVH'.@YY%DT=W%RG]35D>]4)IC46#;BE/A. 
PF#"H-"G@[=$712Q^IC,GLJ!=[;"_!"WX!L/R4.[/6#T!<N1GZV V. B?T$F*#-.D
PEY\$,\4Z!B!S^KWIM-TY/<%G]1^L+X6H I(V(8?\>P5-F;"L\2"(ABP:?(%/[P&3
P4"E1S=]MI*6>& 4GC(+*Z9":.1P!BF1-7))&U,:&Z&G>2<S@%DU-T(X'V- 9&B@G
P92EFIU^Q#EK+B%)AKT\CENC=+L.>5C6(YRP51@;"P(7>&@=^YI4&L,7^'1>H#14V
PIV4MQ*CZ-GQI>O<].K:0?"-P[\9S0<6NT9%"B!?:2LD=\(D<\/P2U3C F!;!Z'TM
PZ;26G##L $'V9K*Y&2['QG9C]\M$S+DJUOM$!^B^I0,&B9G@.=RK6@+I$+&6V8Y[
P$Q\U:@QT%"69'"EH1NCGB,]/>#,PU.^X B0![]H5&!N)0^-,J:99?2_7+:R,P$V 
P 0+.U%0)=MCWIP# L-F[*W"_>G+Q53' ;=-IGQ![6#>45:U4S"F Q'%5!S90T[*2
P[AY7H H4"[;5J]MVK#[W( ,9VI<GV%6)P4Y I.0_FG!,KPFF0Z4D9[(_0,C+Z79F
PY<BPHRD%B@*LRTT*V\Z?SK1[C1X$7$CC7#J53@=$Y!L+96RFZAVK2D;&BA\+_XE4
P28/3((5_@.8;SS6OC;&1QW7TBU/A<!F<PYK,3:>S[Z^46)\4,RC32I:>PF$P3\5#
P%##8 ," #YB1U]OUP8E<O$L2L7RM\T2>S%4PJ_[M@Z,RDU-MVO=':HMXE\QYW,E)
PHT5%Q"9/936"VA9EG4A**KW]GV2QKQ,M%%*-T,/I9 >TI!U$3@[68T_>@!8DZI1?
P+(C%]@O%ZUVKLC2-D&P>VP67:^D*@FWJ+@KY\5USK"2X'I'[O4 7;IO)=4T3]*5C
P9C991*\Q1Y:-PQMG'LUXXQ6^]8WX3*2Z76],> R<1L@ALB$1N)W-DLX2:5I<D^/&
PM="@FKPPJ)WO@X):=[1LXI?X+[N7'DMYYX9,4*\/8UE#R++\3()VAU@=<\KF*\;V
PUO?J:%17[=1,0"^[TNP44#8;>1JX^$_B/72*'.L ?FB:GT==(]<Z&#6$/> J6@6[
PO5%#^3KOCC1#3JX-R*:YSV7Z1Q/^^K W43%G6NA<D[E'TOIP9%O@4MPAQDCIB!-^
PXG2R?B%"Q:#Q:^&Q%:=H&V;\-ZR)WUC1>&?.0CE4FD*\^<T)AHH9EH!)&\+PC(GN
`endprotected128

