// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// File: uvm_dpi_object.svh

`protected128
P5$N&KO=T/45?1<#3ST0#. O,<!__L-0)7P!("+3_W;EL .($:(R@C@(&7^N-W1D:
P]]=B2Q++PP<<),():E"'=6Q]E_W9<+7\J*#Y2%D1@=KUQS70PC$WL*;[G4-GT"(L
PD'H!D3%4.YXSYIWLV(4%RH^JG4E'G9!2_NEU@2D 4&.582Q3([7+["GQ5N=Q D_.
PR=;R&=6$R4Z'Q%Q'-O6KUBR?7? DLB_:]62F?1$PDZVL& <OI@<$)&(Z(U3*8CS1
P4U<=,34KA?ZOVRR%]Z=NE,=EQ#%9T:."_):J@4?O\@TF!9JS.!-EE9M6<1:S&PI;
PK5@WK%W7<Y=!L4+> '1(@9W14'>DW"#*0%*>'&7S"&; WG4)*DA^5"M/]2U]5!RW
P*C5:7W8D9"9*HJ>2&\?_;SMA/E/CM_OU=L _,9XZJ'[G"V9I#EB6(L705&]6"MFH
P6?M;-((O.4MDMOI7L;+03V1OH,7#(+TQ;%C"A!4C^85> FU67]^:"K'--R^%F]N)
PI7)/:#J(X8DG><&@G;<M-"-&8W AG6,"2L5?G9>-TP91J4,/R8G(]0B3?<\L\J2_
PV>=!38:<CE_C%T7^^QO9RY!ZU41:+9=#GGJ^T[*S;G+J[2;;^823"T&_/D#QGM/L
P%SQ\((<*PB5%(_(U5P,2&G2&ZUHG=GBM;'-M,I%_X[Y&ESJP/NV.=@E9 XY&0+'3
PA8@M;F@4_X(#-K6DMIZF\?T).B(=P 33JJG3O$!B3A56OX2>2,IQQ\6TC3WC@F>[
PR#D\!/8BMH@!XV]ERSX\NDDG3JHIB=^&G-U\:8ZVO*4.(,60UT"D03'IDM00^^%7
P+^ENP@VDR,0 $/U$*N$HEX_#YJ/\9XQE'J:#:?T7;AW??KR8-.>1!O/_Y1,4EDTI
P^O[@(WK'?)>GD\;YHJ+[L?0J@2X</]*CZ;-1]K3F0?XYQ90A0MN$/]-*&LR;<HVL
PJGSIKCU)9\OLCLQ9I?V%"#WG#<D<J2!+GX3FQF&/LC/!*$#1UJAK9:-6 BI%QVK#
PK$@J$)Z<T@]"JWB1YH,/LWEA;\,WK!F.1?* $OLV!:=?!3)'LJNY$.G[B<+A\OI:
P+<EH;03!Y1Q.2HB0?0?35.HV8)Y404$P#\(]1X?G]M7QC,OE+[@J^IBC :/@;EHO
P.DMV.<XL5-00.%LL*&FEL%F#5$W-'@8N0'-<_Y+5 8S M/@0N,C?1BO.AE>9BK,Y
PKL:_K=;]]@D N*@.)$Z&)2-R\B=Y)V4)#&P5C"!1XCZ&1R,%F(64"B)T6^X]&@>:
P]TAVQ!"ES1CGE F(C^0#.?D ^Z-@[5N.EYA'RSEO"@-12*C&A&4K6 U5AB?Z<VY3
P!)CPDXN_;E:=@0Q8MJ:RNMK25^7-OIW^7G36D!TACA" @VE=5#;/KL&Z8 "^EH9#
PM1Q,WY8$FP%E.QXILE'180/R T%!C?2,D30G>BUZD&*_Y+$5"5T6BBB,_SA"&5\W
`endprotected128

