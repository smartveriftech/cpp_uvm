// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
P(_+7YB?09[2=*GW'59T@V_NI*3!/&2['0Y RUY N;>B#$WGGU:7A+=DN4^1\YWN@
PF)7]+GR1*=")CN< 7XAC:H)HG&$AFQ4N/";<FR<$];<)L-@JM6)K3)BL4-E46#3A
PMD6=0WCA=+T /<A*XJ-ES?/-BI9O0C-E\)Q$<U]3X]%E :%;U6T%.%8M@"X>XW0M
PV C,G(9V5&90,?<@;?LAFV",]KM$F1*8LH&U-"Q;#:@^";0R!O=)A7A?C]BH^D@Q
PW<TOJ4!4B@%NBSL>G#P,?Q56GDK-?(5UV'<XJVB#AB&Q5D8OC'-@@TP&BQFKQ(:)
P!TTOW%.8G)&Q'SJ^#@L)<<*^DW2+D$!=&\:4]X+H:ZVABYG*%-ZJ>SYJ%A53G1_P
PGTRV=$E@*Q-'^*KWT5%6#Q3A_WJ#9FQ?6X3)EE>,5/4$.1V;&76U0[<;.GH:<ED<
P\Z&W7##S<1R(A*T5F<,;O<X 7*^3GOZ1/,T6T3(W;R8L<6?G8,ICXQXM.>?\_KPR
PTQME&+9Q3;?L8WCO[9QM\L7*QN!?#65%TPWZ@^F 7U/:%\Z!YUH@=8+-D.)'C&34
P%;6[[W..# 03]VUY.8*A8[ICG=PBWR$M>26Y>GKMBM+Y+V,&5R?K^.C<IX)*C: ?
P!_D39/_7/D8G$[,%,Q-<".8?T!^_;$P^D^QJ^IS^7&%%Q4^$BB7AY9_PKO\^7DPP
P&O[I%88N34'Z(LOH<0'PO\$6 8@./;0-SC#TF7T[X5Z24ZW0EJKA,KN3W S5>N)W
PJX4'D![']:T](G,45.+K8^,LYY-L&&KN31%W-U&NWR=-DZ@25!OQ&R28*C6K/<B<
PSD7RAM(I)H*G0JZ-KQ4TV,*\X3E 6?4P((;/=69-[Z#+)OY\F7Q,J1,."^')?$2F
P4# ?;8W 6AGM2X/7Q_.PT"(;J[[MA"<9IEHRCJ2!_>:QPR#\^^AW=D5RS7*7@R*R
P:9G-6N)E .SR> UZ"Y!G"27=WOU[>#;8-L?)JNNC%T[&=D'!8"^@" M19>=P?8ES
PX#T5KW$!5.Q]TE4.]#X8JX'#QDUB\]1^,YUFV.X(EK;^B0F=R_OR81 R!G'*V=@"
PG3H%5\+FV[>BP[4(@2W6OWLXM%H;O8U<^1 A2V==U40LQI=Y/L\AM?P9>S=7V_QS
P1AFMV; SFCY"\N3D,6&2Z&NPPA'+>-RI+'^-E"*4.2V6<UQX*4P=0,C,T^1^L^+3
P'OT=1VCH39*(_-):QT)7M1YBY=H$.,D"]:=[=!6GYX/IQ8VN )>(1+C#Y8UV.YV]
P&):L=ICNAPV3#0]20Q/B:=Y,[J""P/@,7YXGI'1$QN#>%3VQ,76#E\IFLU\'N'.R
P1VW/[[L,)1A-\E@.1+(H,D0DKZME%W&Z(&L+ =@^>J]E8&,3YL"9@8:R  US)$ER
P4N'[M[4^NS368#?^P)?_'#>]K1W5,Q2VL;]JMYB#LSUQOHVR-0,LD9Y#R,6HSM9?
P_WW\QVUR4Q!=,^4?GC3_0.GV>M>;3VW9Z0O,Q12_:NE5Z 89TS/2B?!KRTK7&4G6
P\\?LJUVL0RZ@K#^3S;H!R: XJ.<K72F>Y]&R'V%[>\#,F,7Q/=+R "WM? 95C'BD
PA2VFST=4VM<I\U;15^]4M05M0Y!.\63(JC9.%QI:V7]A,&F.R(/5UL5J+K/!"[T@
P^6?A W9GLI%DH_&(S9.A0&35'A-<H.3B@>=-2,_4F%U+,R:B%4\@'J8T]5/8%[P/
P%[[N1/==8+Y[.&:@Q](<%E)SA2%0' %D8<CRY-FH)J/BD;SO2KUFM81%-^@C>8)=
P"].T5G^?Z1D:= M;Z6MM;/4ICDJL5G(/IMVOK>-.R<IR.V_C63-R'WPEMX;(18;V
P>I"AJ!GX?0QZF2O@&@8Q?R13377-CD;'O[V'UFC0;4QO@_82+6IYXYRNHSLA#%A-
PT]Q;^/!Y!IL*'P-.AN88+=)'HSYTL;2,H<@E>?4]0FUQ8R>0(#X-+K[.N[VN4B"0
P/\D*@SI(/K4DID^8&9 /'I&5F6F;'[M@_#9H\\J=A73OH4I-CVY4G:S<$MOD8@6K
P6/E^USV!S?3(D$W*-:U'%S$_TI";@KUDN0<1V#BV+;2I&#*VX#!$GV<4WDS^S]\M
P$POA 'K@>_)JBND-H:K869UPFU7E=_D+KI4OQI/]:LS#/OY[(K 3/0SM/@;TL\O,
P0*?!:\<8%H[TC'N+QG7[LO[R((@$K+LR-;!VH52?9<Q\WG((%H+5H5GH4I4L[A B
P<I3?08U#571<JECJ[.FN/RIAMW@2AW9XQ_&3B)4-FN-L]Y2@:+KZR>53$-(L!3^G
PV^4?2*5,L'N*6 6PY7PV%#]1^F*_TCAZM??DF7_MM,T"6H<*+,M\SF8*_=8 ."&Q
PI.;$5YG";EQ9WU_G!BJ 3U!BB<1P@8I8AM_]6#!.K&CY,;*#?(G&/,2O?E=FRW/G
PP[0A$5OI2CPO;PR13A$!V:& /:![<Y9.YT:,P0:C'15VS:Q%JM>?T)V1'<2,42M\
PZI*)#P?9G+HVZ]6:#[>*P7'N14-DYV?L)UHXUH/91D8B9W,K0W"%N)0>=/F@ZS)U
PQFTLZWJOT_[05[/@X[$PS%@BFH CM0[O2BJ(^?ME4_6\QMNJ!8.S&P-+7K@VFCH)
PRIC?[DR8(R/K'P^KN_#B1-*#9C,3G67[*(?-M4<L4-;H+3V<GDA?N1:K"5QM'B2-
P3S"?<HL[\BN=A;;G@Z@+#P7N9WFCA]IF;N!/4#OE<KS,EBXO;.W(F!;M7*M-DENA
PWB5"P<WM2SRJ=.I95>(&'L;9);[IT/'W\TOK,-WJQ>;!0'9)^6P=1K+W3/N(=_ZL
P?-<\V":T&) HD<1N-5@>R,1\^OL'^17&[J@;_P-IT(.UXI;RS[@97=WDXQ@WI/@"
P@I+M\9@BUW:G4HKUFZ$.U3]VJV)N8LRJ48YN*H.)H8Q1+\!4K1$Z7,WL>?FOX;^T
P']:[(N5H/;>H';%,/Z_P)EM:FMT.,TBRE5H9;QJNIACHKCQG[39AF?Z'^1[(OBMO
P4Y<U!DCM'-BBUH.=#H:@-MS+OTNR 3]:*?(!^U5F9286(?5]Q#ZG*Q;(K $(M65H
P\@SF9_=I0-OE6 XO 0ARU1FS39&3X2R@!7JO/Z2UM+1.^J8LU(S<L&9)#C6RKXW=
P0= C$^!CF*!!+A2:TC4:<QRUS!@/YD>% /13DCO,KH2;%HFGUC'*RLXK^"5[PF#Z
P#G:'1]?G&@/@42-P'6Y/  ,QIE(1V>\ OVE_T M=U6A&[Z6C*FTP6?ZN;F4)K/<J
P==GU1<9N*K8W7%7D-;+$>A;F/E'XDL&O?7W&@J#SF*NC*IL41\;4'/*1 U'=VY\<
PFQ!PN^N8STB8Z+.L<Z@T;)0&\E6DE98 \N.')E-378TQKS%D>..6]^IG**/T=+!6
P#)_+@:G+#HEU!NHZX'S$$;>OVF\XW>;Y2'=[= =M1HAV1L")^54N8+ZY=H,AE?\.
P<X*)/D!WM9RE**^*<>\U;OQEB8';&S<;11D/046[+*\BZ/_@/VG_*6QZ&7C%Q_SN
PEVO3<<5&/USLB*O- $=N7]+_>$\07>C-RR I+X:UICI\$Z/*2VU5Q#*;U*K.+6-P
P5:'.E#ZOO]]8B@[T17_48G(":MO[]E3TCG2T[ZT^"[?5N$OMP409 YZ"&^,8)B4U
P$5>_W+0H$D)#-R7" ;%SSY CJVX4Z-XZD*$*EHQ+ZW[FAI<FB.6K2L+.7["\6=(Y
P6J5[S_A&U,>4Q?$$G- %=*_9&S_\L?$AGR$@1YU'V_[G#A&BE^ W2ZJJP&]\,T5C
P?@9//T8TG>/DAP.B/JP:I KJ=6!-S DKFL."HMB>N) GPW )00/CKZ^!)K= Y0.=
P;SGUF=:7YR0C'W(=MILW@_J>O0P[K )>+.Z XH(;7LPTZ1&>5LB[QT) YUJGV8+*
PU3@Q*D&*K$#4Q=GGYV/%!58)U$@;#6B9 ("=6@CN0.+UGM<C<IRK\P_ENC0RXK:G
PK5>#.,FC5AHH75:ZWG<KH_S]#025\U#R/X'2JFZK2*5)5D<5\0 VCJD-X#W6,FW^
PV\LF(KSOY!5L!Y.*O$T!S=-0LZK)U'OQ-^P!3MLOB\,<+'N8R35<_*7KU[:J*HW.
P2,2RR]QZ4<]&6G+1>R$DJ>?98""WBVO@6M/7!USJ1C$#^K??6U^5 ['P%?U#R7Z)
PI7)@_@6! 8:JD@)B6F(;^=D$Y_&N/J:HF;[X,1FNZ[,8M5?U#P%DL3ZH/H\8_ZVA
PK-8M3B:3QD0F?)P+/P<P?)1$5.5T\SX4E97. [0R2!5K/88VL2JST#1T"XXX%(*8
PAS]%<<L[SL+G^^ZX4.N!NB\O]$_M1= M.9HJYR5^T/;9XPC@OF+6(^#M$N9&GVR#
P0I1-5S@!4%9?K*#LI)=-BPQJ?6\F"FOT%$\(A Y(RQ0??\GJ/.5%>E/Y^S2JMEW>
PI;D'=ZW?-!4;HQP2Q'F[3XJEI7#J5-J2&<9/:LX\9+,']I[TS@L/R^MER.5Q(1'9
P+/*@KO+@_U;MJ2W&][D&;.N)+#J]Y-@6[R^>#G2#G ?<H!TCQZ#H.F[+*QW2?)_-
PS"-(#I@Z\8F9V:XX<<7.GGVF<DEMK$LVX-7*H>P=-4=49O#3CZZ="A!5;XB$('Y"
PB++=6U4;4<.A&O%SCP *:FWIFD>,-)[Y[RH<7!/.Y[Q8U/D:\H8IP[ P@&ZFA@ -
P&T*P?WX4DTM&+R9Z@GQ>(]#U'_L_TCRNI89$NR_XAI%INK9CW(-Z#%>$5>B&&XBK
P\BC%A$45Z)'((.8R9"$9<H:V?2NU()]C7)Q0@&XHM Q5VS+R4F1)V>N<CH>HC<<E
P@O\FPWV(_N>>5XY+712CTY1 *D_E'B?BPD*N]K3-X)5P@A4-]K%:1STR*O?3K\Z0
P\?'3@=J;IBYC4MR$=[)6)F?*91$"K_Z*V)0[D)D\@P#RV'"\!&94 H6^S$]C+?H=
PF*<H5:WK;(NF0]=EY@>@ JNL[WX;5TUNHU$]5AXSL.'_MTG7)J#7#=T]SQ7QM#'G
P1SEM(X%>POFG>SSW).>A:C&LA;MIPT+([$U!81[+YCKOP(%5.^)#53^;I'3Z:26=
`endprotected128

