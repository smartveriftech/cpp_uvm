// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Guard to prevent multiple inclusions
`protected128
PJ#U?;>_1HTL+FZ$,/VA:5V$ 1AD9UP<B 8@>42H6(>A&,BQ10)99A1J["_;3-I/\
P=#+?>IT%>?(>L($.!XKTS%1/5:-7,B>/2O!;A(B9Q-7ERK?+$%&5M,V=#C9AONV6
PKD6+UV7JB-),8W1=HU"81=R$ER/FJPUJ01(DZD!F,_9D]2P_5B=Q*>:F&HVO+M1;
`endprotected128
`include "uvm_macros.svh"
`protected128
PGXB<9?F8-<'W7!G.$8/M0)MS[9^DK$-9,3NF'F\$J?%QTVG$W:2#CJ0#SJQ%(K+E
PDKZ2(ZGARSX7QRJ]3+(EEN4Z^NC> Q(.:6*FR M[,#TJK!%RD^$O#>Q;2/A37UM\
`endprotected128
`include "macros/uvm_dpi_macros.svh"
`protected128
PJ1YWBU,0,@1NUY2B._V.>4B'C)F(;F^:,#V:4JS>"YP8U@0FTBO"<E'^&YM>!?ZC
P9?X+8R'( YY[%JTJ*1XGM/VJ]+B2OK[G[Q9-$>F'"D7BGMZR$&Q":((?D":6FF8P
P!UKBK'<K]'"(#@Y$NFPCY)ZZ>,'8PKO+FYK6W,<=UKE**G8505L_70V24*8KEO_#
`endprotected128
`include "base/uvm_globals_dpi.svh"
`protected128
P[:VW*+W<=FEM70RLT>$E/B[1+P<$='G4Z6P"W*4^K:@/9B!=62R00\4[/PMY[R1$
P%3Y[9\V;[32[";FW'([]T\BW%9%G$CF@P3)4R6PW(=%3-O1)D_-,4WRG-]3V9^<3
`endprotected128
`include "base/uvm_dpi_defines.svh"
`protected128
P_\JF.C],1TQ2GL._&?',(1^L\LL'V9 R387+2XR?YAO?I3/59355((BXNJS(/'QT
PBG::;: T,@+8G8IF07;V6'%@Q.D7IHJL2=4)MMJV4D)=SVB[M9+=)NC"& 24GAF"
`endprotected128
`include "base/uvm_dpi_sync.svh"
`protected128
P+9\K*[Y>D/X;)%L.^:ZI$V!C:?5<ELN%->.IN/X,N#AQ+:MSS6S./LG@[<,I99G*
P<SQ^_Q?'F?57;$]:TLA(<JA/'"U33R%&A]!!D0GM(7_[ !\ZHYPS/!K(G$YHA<.B
`endprotected128
`include "base/uvm_dpi_root.svh"
`protected128
P.M^<20#A^-</%4Y:JU)W:-3>$/Q[D1>#^S9'*.ASH0T-B;JHG@A$>K3%YHC)R2QU
PLK 5V=VX>W KZ99NJU!C5U0+USDP0WFARL(2?[^U*BL,'X1D\%<U54UF>GU$^Z7M
`endprotected128
`include "base/uvm_dpi_component.svh"
`protected128
P]_FY7'2>-OHCBT ^#3A7*OX7XGF4FRJQ)K#0E28I%E? ,1VGLJS"=%WGJO]:(@'6
P-MS;EJ) U.'&AJ]U,R&RN=)LQQT/L=G.4@@R\\QB/TTFC,E0G$=AA)#K,$'!G?7K
`endprotected128
`include "base/uvm_dpi_helper.svh"
`protected128
PG&#['+_#9D#DE#PY@3+I,!_U"?WJTY39O2"+L]C";!T-Z; HSUUT\2)Y]E6,_F%3
PQMB\B*(P:0,*!&L"PYJ#.O])A.M3K'_GW#0Q(X%]N!W>>:N6-/)>^5&\;@(9AFC'
`endprotected128
`include "base/uvm_dpi_object.svh"
`protected128
P+J"1-S#K(L;)-]/Z)MEY<.)H\ZOY557_4E4G,D6N<-Y5H1[OB[O:<P/+%T=PJ &Q
P@!W5 ,4?1>Q*@A-UPPXWE4G1^23$H/3T:38\&D=1E;)M=VQQ<1$*75JQF$$#!8#)
`endprotected128
`include "base/uvm_dpi_seq_item.svh"
`protected128
PA+0/_DL\M&V>XA[P'WX'I"JMC10"I\]U6.Q59QAY4J7\)N68-0M6^GR.9,K3EV7 
P7P=5E04E?JE/O0?W^JSM/*&Q'^2^^O$@,PP?<JTP5Y'MXW;/$)JT912@^'#'589>
P]J<;P;T^GE<-%<TJW:/QJ1Z[,Q5Y"ME +3U^X$</WAKB.&81-H_B/'42=%'RS_2 
`endprotected128

