// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// File: uvm_dpi_object.svh

`protected128
PRRP$?*/2"RO+LU^?0CQETA9F>=6S*\XTE<5+%O1/;E[,X6])M_VY,6]J^$>NZ'E,
P@^3!Y:D"JU>QN]K\X!+E# GH_\99X"=("]CVD],ED^&8YY)W?A&2JV^*X)N3EF'!
PS\'I*00GZ--AX6Q?90K+U.Z#EK79=.+1!RT6MT#_&B5&T6%R)X&#-7S!V_,;ZHN[
P'V&PN<P_Y4&VZBPBKE8O0UKSK=;XV]S37]X&=E$Z;Y=B1WW]A"C@<BM'5\NGJ[!M
P1!,GD2"D99XKZ]5.74Z>'^6/3.B29?>:;F(&Q"+:>L8DA(\=-=0!MH!#\*TQ;65(
P(<3>K&WE$1^(76YUZ"N,Q]S>J]A&[<!^WJL4KNW0-QU;8[Y<P-W;R:G%UC7+_+8 
P;P.&E 'SJ8R-+&_*OC(EDI/M+))U\$>?,2TRR;>C<)';U"SL8LG/KIR@6,S8#2=,
PPTT!:,A2?_[SQ)S#+E6*OU(Z)Z+;80KY*\)<]NF]!_OZ3BUE^^>C?5XWC'ILMC57
P4*O^*HSN/OJ1HAY="08T$):6>U6"G&#-L+LY-SJ_,N<5C+@<3[-0?/ 5LT$^Y]QJ
PT7RT<TTG/Y&5/4G3+["N"P0,E(+='3 W#.^MMW*CW@ =PC<S8F3Q)Z+\J2<3A=/E
PFJI W&L]Q1C.M(^YL+2=9\!7*WZ+<>0/&54;RL((33XH&/^G[ZE<1B]L"G3RU;]*
PV .TQ2[T")NU98E;3&P: N:9Y*9"QAZ^,5O<Y<XOS@/^/W20>./YJ.I)&P]H_+#$
P (3QQ>/=0 F0 QSP9G 1C[;-D?@](P50>\S@_?0I?#@S"U4?'!2)UFN[2"]YS6C8
P-Z.)E]=%2D]]('4>^YT:'(TN2%2/*MJ+MLI1B X192&E@ 7_A*50F,87<57LU#BI
P/( H+.N757SADQ6?J:=LO\ ]OB$0/OH2PS5;C#G+:(43D2,!?X6K?=26S+\,'#- 
P_T?<6VZ8THMB>N-=QBY7)94J*%V==*@VJB5O=_,&R &SL&!),<-'J>ZS>O0'G,6Q
P[NRYN@]P6W=7O;J3.8<F,M] Z6K*@=7/!Z.87B);9K*/J*]X,<JM\JT^96_$$ *@
P-K"__'V=Z6 ?.=Y&@R$MK6)L;=%"QDT( GF"M?U)(+%OH%Z>:$V42QU5"3)[7N@.
PYM7J)RU0FM5W?^*S+0-I:7')5B35'PX5UPHB(IZ[**VKQHD[MP=L,UV7XJ)Y2=6)
PT5WYR(]&[6Z79DMKK:8F+_!LKFK+-]*4]0'BW!4K)C'(C]$5FSDG][,[3@B7D=,R
P?WQA^_1B:P'Z!N%H2WK ,!^OMZ)24$/R%I<=*AGIW*+P531:B5O -@-F] SE+@GG
PXJH \=7NB;]&':I$01K(A3M?Y:<<#<QSK%X) K^9V]P%5YW>@!,[D1H':) BRCEN
P2&[B^KA%NOW !^,[:QV@*8,6=E,^I-\,_'(TU2#K20DFN0*D,N7U[5O=80<(01?O
`endprotected128

