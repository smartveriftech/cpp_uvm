// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// File: uvm_dpi_common_defines.svh

`protected128
P.[\VT!N"@Q&4K$%:.LUKU3VKNB$1-E9YJ#8.<\Y>KX@<+K$Q>6QUV@S#U.ML$^ZD
P0LR9_+4N@-.\.+60%R=!V1KSQ90*!G?;N=T12\ZA95:DC!.Y:KU\D9V65QL$J=?G
P"2WL<K/ETB66I0X9L-ZS28K:!%,I[F/9R8QZ*7X>D+<F/ZKJ=3W'Q]W(5Y6D)&)4
PD0V3J#V-@A9Z"/L;KW\"I!:<QN@=3XJ2TW5@-PYUX"YGY0'[Z=DCH_ [MN.B'SZ;
PSBH':7MJ5S^['Z8,AH.U3"9]F>%O([QQ0JAA8& \N&#%)-92$'#RQ*_XE7MSR&]F
PNCOM/A-=\%AC9W8JHFU<-P"21(%20*0Q>KZ&O!''SD&9B<J$X)WVUE;@9L4VF H?
P6"-+OW]_.JEUBN='B.K@:BC/<[4P.<5G_Q2?=UY^L__BM!4G8^-Y.C"W&C7D>"'6
PCP!CE":!$'<0W-+GC@0?F11H\*$,CI^7JFP(1TG6)_N&PC@??22+ZVQG7QTL*.55
P$V::Q3"EV@IQSUQM3@6W>;L':T*702-4.@<>S#^B;\*D<0Y0>5%)X-9O3-U>>X<V
PMLF>POA(UVU_09[+$19?(4D:Q:/-FB"O6BOP"[;=4T&\8[?F"BJ,JJI31AO@N:\F
PL7JP()=P>(WF^T+D56+B];A>GEF[-X>'XZXY:2Z&J0[C6G%4'TD#]$DAE8O+KH]T
PH*P2+)L,V @:A!LLH3$_SJ^;0H<\G;9)3E5>\)/\4D;D&$T9\<+$%;(HR(T M;6Y
P^Q8(1_8,EI76NJC ,[65[?%?'7*RL2C$_7G\8+)@D?K.2@8<)BIBG"KLE_*425I8
PGJ;O%#:N T>MUGE/$<,HM5;.]UFR+O1O2[:2N\:<N05G!5A?G@]_.7:C(_!PA%8[
PF8VWQ<P6 AF-B8%-6'*#07>;PL4Q=T6^6'^J845.*[A026'<KT11X??D@"/;4WB&
P0GB9%LA^PZQP08+K-E#,1Q#,G@H52#_J5FO4MSU=TL)7]5 Q5)-A#E4(D$O^ZP)G
PJXLNH[]WR>D9Q,'1?S(KY;_WNE(KN:I5;ZCA7D6X/)YOH:@F<O(43L>50;?L@[JJ
PW]1:8+@2$+2E\ $2A\G!V%G,+OR">X>UN54G-K'<083,T]I%"3)OL*Z5<*(A4=*,
P.(,K=8TUV*P.U/IA.7>V=:Q9C*%=R!"LD;A+J/N-KL!Q"L#4^ 991A96Z2:KP$WD
P2<M"<N\?AEE[$.R]4[V-M^V3:#4^'-U572]G,<M]7CD ?18CA-F4_LVTHW%=X^^]
P:'+1Q(Y@1\:="UTW;:"O74K3WZ9+&>&"QPGS<F4XT5V3A;H]K\F^.?>IK*OEGB"#
PWXZ0BW:L(ZOE^:^H0J,;603@SB><BRM$;!2$(R. 2 #<&O+3__;O1CY! L^3O>"T
PS(0([GB'UM:>.FD#7_'8% Y>$@$JH1NY_;D(*>K>GN>A:WI7S)2=6[4)B^_CGM5_
PQLXW>>W'[*<=AT:XFCG\I[14%I[HP@O&_Y*^:4Q+7@/>_F<"9A!!4'\+1-%5!%G!
PA!]4AWUA,H=[7+\FH@3H&\0J]DN454GGXYLPP7+!PMBEVN>C,JN^(,\#.2LD[:Y)
PY' K,:$&']2E5)T<>-<S/:TBU^.B XDN1L)AYX7ANRT0:EJN7F1>]40WO +3' 10
PPH[L-M,@CA/ZY!N.4WRB%;:Z5W#_^PTMR':GBX;GAZM%+";L"*I6U0\[+KPU?*4:
P)_CR&%@I+/USU-,@)NP?_0;^BS<29&C:'T!7E^Z9MWC1=,C5Y,C<^Y2G(? 0GZU]
P*2?0^;A&%RQ8B+V.'OB(KO8!)_Q[>[D8V"@/G%1F,P/_W5C?!FO!1!D5!F498$Z1
PN6/+.S,H>JCXB32'W0QDY'S!!+4Q1471-J3V;F:W/FB=S)K&D4V.Q#,V\2+,L1!P
P0* T'A0CA/R$O7U2^9?#'QA<@/F&!$,8?V@;/YD@H";"G09\&%0EJ"N]GO;^(5EN
P4G^V4L:80O3>W^.Q\L!<> 5M2$T'UQDV96;X6'[T!OUH&&BORTP9NHE [3/M>6KX
PVCUQE(S96^'5\RDY-R[%U[5E:!SRP@;18YB^)#1]X:!,YR%I=5&6-JTBHX:@]D%2
PKXCWI:*F'T:33!T*NGRULFTNF!U#O+CU]_RQN.^E:?$3^7&MCUS@ZRFAAP_WH!?)
PEGF^F:>Y=X^UFV1)JI^NB!V!N=_Q XQY*LAB4YFOR_XKB5&1$_,R(P+ Z+S\RGM7
PCM,W&VWBZ)=426852WZL8$C9D7^[T$*R3E.L'@'3?W0P!1:!!@PD&UAKAJ$D=WM]
PII77G)$"RP\H9.Z\$\U5BN60K,#@>I8>:.E)/^0',RZ*2K'-"DH3!/:!B!2E#38A
P(86@6G[GJGG!MN::KYYF;0W()W4,'0QKYI$W?>22>W.3U^E_)ZUM+4^%)BS7/HM)
PKC3AVS,XO*IW;OG%J M?!H4.Y&!"AE:2'O"*3>(RJ)E7-XX$Y&+#A)TO5KC0 G2.
P:C]]EM1PT8^9IX=8R_'=-ZW];U49V'_1DOPK$J^[:/XI#49'C;A\=F,\_=*+=5^4
P[GP'AVFY ]Z48T94#D ZRL_LY16#[PC:OIW)4#*K!LJ=6M<GX)I>91=&P0,')U10
P,+ZV%_N<XL0VJ[PYSN!]%BQ @]C-^9(A\- KBY@Z6:!9QZK@+6,(Z=SH*AC&*#'L
P<2F,J$(O\X!120\%-)IGJ%"#O&Z_P*)Q)6(NXL'JQ-#8_+HCBE 8'ELT?+> _,U"
P)B;1&^;51V[.DU!%RGT3$/$;5E?3G8N^ON9@=D/Y$%0OA69IG^V_C=*Z8*^K<5O;
P3#S@@JD,G(D2VOI1V6"D>N;_%?K-S@38GKK'$"Y2UU]PVWNC9_5A#VB71@3YHT#]
P69$RMTT#<DMI%E>.%6;9>Z,Z1KDDTJ5MW7D5)"R(U16 L] Z[21BP88MX;5:_RA:
P8 ^JU>O=!85>G/$$T@R/^NA"//ZGCN&Y_6M<D"DJ,7<J)CMQ.!!ZA0-LFDR?._I!
PG 12L5\$"RD!W)GP?C@600W/:F7@2C0!WZ;AD0,+6G]+M3RE;)8LIAN5$$Z3WJK'
PK1+@[?,X'-7B$"+\N!>U 1Y.5^4J82/(&6(4M(6 7!;>U6%:/UF\HLMVY658(M9#
PK).5(9=AYV1U6F^H#.+^A/K.^/N#A]R/CL)P1>E.'.M90!F47[QGC-7US:W<D+)L
PM;LB)&@<EUI_O66:GN<I+A<ZZ;+9I'<3]K1@OU)/F=5I-E:2B7#>]C=4)ZJ3RSO;
P''G9", SY!?1__96HZ)TX6WXSY?E;=1Z,"'QW=!C:ZM6)8*D0(G9KUH".?"UBD#X
PS FL2NPGYWK+16'.!KCDK*>_$:?O8HM8R.O6-8XA?7B,L'!Q >LNZV+]'@U4U?F4
PILW";8[&>+E-[G25R'QUL:UMZ=A/SKO<VDMD;;&4IS(D#\WCI09:/NFWL63L$0BD
PJK=X'V6>J^>FKK7=>L]S 3/9>WX$!S?*BG8GSG\]J9*]XBKR%OPW;NA0A&/_0(KP
P@KB'=D]]#;$1-.7OWU,U_*B^B"D$M7KY0@'=5UPT1CS@A00PFATY&CX* :L&O] C
PBU-G!@41') U),/B"Z7M6ONC9XN.=)>-0*<;A/WFSN,#NJDFTC_XU737QS;7- @J
POV&<ZQ?@8\^6"?WZG6@O_5A'&('^5WVB'<)9[08(N067=O-#CRYARN4QQ69D22D-
P+(+@:09CB@IN*U2 J'U )1.N8V=QTKI]R278"'H]"O^6A[6S(V[]4!X">J[&%X!T
P)6K+:<^*ED5IZ_M\?\1Y\JO-1;%]E-><OE9X6S=F/;%5VZ!UG. 6L"OO=\<B'8PJ
P_&_U*$&X_]4,5Z&+\%$O(MZ0M7S"/0@S,$50+_C.O2U(C+(DV97#;F.DU)_AW@(3
P!,#>3=;M2'K0R47=DW[,L-6,=MH92-#CSRBV>(*C:WR*/AK,+4:O)YRO+P&VM&0W
P7>0)TOD<O[$-FJ_E%8($/T"&_^7,-ZM!!2![I0\^"0AY_4.SAN\,S\207XE[M?7"
PA%@^6VL,,537V5CZU!D41*A#PK.T\0?7R\]Y?M8T@&/.M'D"7LQ"EXEG%U:E;NF*
P@\'6@,9!+8P6$7\KBCZ;CVSXY<&Z2?8'\W0/2C\_/';E)8 4>#2Y;HPM.P71:>]3
P$U%X4\ !*<^]+RZZ'C6&)&_5;C?C#.IO9=^DQH,\5XVAVHX1:%$-D\"90?U,IRQ4
`endprotected128

