// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
P3ZUQ,G>U/CM")P:05,);=<=K]P7Z6MV(^O]UU/!K,Z3C/_3%M40:?_W9A=:BRNS3
P!^9!EP!ZT).)]S<?>UD,KHWJ:I_ZF9N;;<)=^&LK< T)YUT@T#>%+8T&0;8/$04U
P[:5*N4:*)!E;-;2.E-38G.))&HTD^/\=<CFV(\^J99M#JR(T@%.8&A9)1_V]/W2N
PB6,OX%,.82L76W/QY.$CJAC'1L=**JN1U)FIJK@\1$N"TATK-OP,-WEES\Y*? !E
P"&Q'QC"8F,Q\225.CHL99X@E9 @>'&(.0D?C4JSQ!TE;)C1#O]FMT.E02^;:3Q\I
P+$+^/>5PLF>I#D920?Q2C%^2GZUICLEJM$$"P.PH96FSG""V8[7-N6(NK#L6_ ??
PA[&2X?35EHO-:+T34OH%0+(34;B.'S7&J#U+B(NO?6<IV^9[W@E.[)^P:/P>DI+D
P SQD\@*=DRUW@[CBQ>(G!6C31Z8E]\8*F&A_$4NF^%!]D<GUW4F6-1G!174:H%('
PPD<T))G'0=G><\C"OEO+$U&)%XZ3:AC&*^M8<1 'X>69J7W?F4)H>'P?BOJ=%X4=
P<@U%;#:DF5-[%0>@%H31ES4FW49GM3L[L9.4AFM-:2D?:4,E2ZK?AH+@7'B,KAI!
PZ]OGUTDIR^KXMB4N56F2W+#C-@P?OU5)/[XI:W%'4HC+V+%+.5;:9@B;7+1&#?^C
P.H%[F3),FL9@QXE[J4Z,X44X12-8?205.^_P>')EU:YI8N0F[+2.":"5HVA*[AX,
P@J];%CM4'SW0G$7-*6GTVAL%MQ(,)4:)Z7.9YCZ-3CN?SF4EODO)$D2O("QDH>F"
PY W!'LSOV/B>(6)!(=,)1F^ D9AS(1<SF!>=83; _NX9=JL@9982:K/\OCD57,]3
P#[V@2W,H68W?"]G3?L3F5IK[!(-"X([NHD@N-"#!(#)N7 MI(2>0WX^$:,/!:I>%
P>-FMBT#A]40U*8!,3GK\WT P0$[Y[I!<>&[URXAC.S82UG/2*O&7\[C2O07^PRLT
PJQ8P-=$R.6.73\6#K;3T2'E)41<*,OA2YOHGO[[NC?;SL)S^:>T_CR=OO$,RC7 R
P3 86%JEB]L,@J[@4R?'(OPK>TPX#6OL*K1IX==^89TLW+9P19:0"0GR:0G=,I%9@
P;#:'#9V+MHX[RNY% )1.ZN^5<5?:^I6)D)K*$@D.!XB1$VZ3Z^8/[S 7NP7-XOT!
PJ=?#HHJ$UKN?$+4PRN.)NX;4U/@<BQ1I$HW_6;:.(EY8>]BO8GO!AV4\_/ 1DR0&
PY9KS:_$:ZA3>I/'SM9K(*F' ;YUU<_JDS>4_0.1(%1C+/ET9M#5G:RCW*ZAL6=:U
PP?'AAE>(^&)PF6C!69A;Q4]ZQ@"J#U;+ZFME!,D+/(\ZA4+OF:FEX+:0"N>MGCFH
PO +,,$N RGXB3RKY<_I(^(NA U9;&GF(EV@+E]>%OW^]^6N0RXP!J6_[YZN2'55[
PIF&),P]OCKZGGU0&VK.MV@\KIMK%ZP5/^YS"02'S<SQ/=G1+"^V[0R<5M#@-M]%+
`endprotected128

