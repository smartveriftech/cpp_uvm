// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
P\/(_ 5<1LD6"OG8+"O1.N(%+:^E0O6%Y?!$%PVUKPX@QUG.=V6")/XXRDQ0,'R/:
P_VC^:U,BQ+W4]X6#='?9DZFYJ%1C>!4H"-!F;90)6L1OC&@S=]T/_*FDD5$@SJ>-
PO#NZ\M\8Q$%K+\R(V0A:(U9_(S5O/?).A^)D2(I>+'Z7,)[7'IY0O#>394TKLXJD
PBQ10DYH;@2-B=^:Z3*-9+@ 95VA2B07VU+XZO<O)>D 5J7&")Y5[Q]DM(T54)L"Y
P/S8LI=2-. )S7=I,!X^BP9K5<0T.N]ZF7Y&?\\2GIGVW>[4N5O[D:9PJ<^L@B\<9
PAT#Z$P*MYI,I^]2;1B80X'24HV?\OOMNJ*W>+KZ!^:I<^F-4V\0$,^1DWE+2E!2&
PQ/G/Q!6EA=@0">,"8T#7@-[+'V<,02W0_,B6FEZ('8K'O$42."=60Z6B0L'."G#R
P37>L49!9JS2Z@*#%S97 !R3U78?4 EW/T"SSYB(&3F$CG<HQ,_Z]RNY04#;!HGV;
PUN'#)N:4SRP=+3T.4!_A\]'398T0RC!+>!&.QQ@8W0#:5OM.-B ,?V'>E<A6'87J
P#@O@A@?K+0=LXNZ3:"*H4#:A/ H"(B)5CYE$[ B5E<QHM<GWKE8!($W>N$R#P4,K
P>0?WW;P@+\4L\//E)2>6Y6D=;*VX!7:T1Z96\N\U.DK;^!O#JLK<\=SA;;RB$4A 
PZ:!(UN>HZW6*CT[#O%G_QR0.T];!F#_F@C&<N&+$6_:3HS;>6:X/VQO*QT_4--/#
P"V*"%+,K1CUQO#P5@GLHIU'910N\I[Y @]%1T-Z7%8?A324HZZ"3:*2M.4AIXTQ,
P")O0,QE)^2@,>[$>V#8@"?", 44FAK3+E/6]P95SXN055)$;W5WN2RU?R:98VE5+
PS2KEZ4RL^G8[F]H#(]>>A\DK<D(-"<5%0!?QN"%@.(".6[[#/X#ETIN#((*'W+Z^
P];S]VTJ:^#315'))']B>@'ZY15](2C<PDY]\K+4#5WC!OKE:/7B]CS_S\-7/ R#Z
P!QWWZS/$3/NCM7#1-,,V\/J',/6]65T<0@=C]$U68N=<_CU&:)!PAH"7-1JCIK]S
P1^J\L"Q((&/ I\X+&(T?9-(TEHM'[AK74U7BF;&>(YQZ]HZ9O#&_SL'4?+I1"[)3
P:^7[RGDL7SY^+U.3/^KGZY.<0?Q>T[,AL]K&6Y/9UV18EN_+/[WYN/X/CIS%W0HX
P&>$3W[@FB:5:51 :^/_47R1='RT)$ VN0&$BTZ!)'2R\B-O'^Z@/AOYGKGK^*>W"
P[]873B<F\6PUQ@KWP&6B'C^VDXSQZ3=[6:-^?0:5;ES5U6"KJ+N(!6 !1P+YF1CU
P'VX@\]F-[R_CC/ (PZZ1'&7(<E45XI<?,-;V)SVO+0.@A?$5Z+O\D0RV/FV*^7;K
PK-3<NBO4*OQT27PT=.")5QD0%TZ(F5P6I 7OY=-AA*P0K?)5A5!BQU!BG:?T@<$E
PJXPZI$O[AJR3WU(7XM0TCA31!=#9;. TW&9R*I?7V5, 3W>\=X1,R57M$$YB@]>Y
P2E9I0SY0VW5.,Q4,C1TQ)"FV:/7Q WO"[+N^OP7*J7N"I/91$@5NVP'[W5=*I*^*
P6$O)PFP"$#<A%?HYKWN-Y/V_2'>A<I?FT:M9B,>%_@+HN1PU2A_%$@?:^*0YTRDO
P&L<#6(_!K%GL[4R!WY&H!?44H3+_!+AHJ7@?_4:MZ<T97R\EV&09B+-WPH;S%6VK
PBE)%9D0K)^%%FUIC7-7IP8CQ+0@<:\;LI;'JG@8G]RRDZ)VI;5FJFS.M\3=/A[W-
PWHP,@:%'T,Q(2 V]+Q MG9?,EN9.>R1RQ(YYYQ8=C2]\R]3> 9N0J?P)[O(:?O$W
P91;":W^:TZ]@YU@]H 2TO55G?7RRUQ9+3Y@97/PIPM]3&]]/[K6?LJ7Y*%FW,Y7A
P%MYR3<%?1OX*1+3B(:$M?'=,Z?<I CBQ#F5*(+HVCS'DV#>IF:M*;02^R:Q'MNIR
P'&HX'F>@&(GNL.:=VRX)A&S^Y8"S-]A_$BURPANP*_-%_M7?^:,O17;$;M]NCA?2
P;AK)'^40:I2&H."+Y#!;;/24PW287-"@T_ !S0Z?+1FC\!!Y*!E%T)7VEK"0B,OT
PW;&%P5!&P[R)ZN2YU>5K3;A0?14"5?EA/+L3AU9^-UXHDHSX/ATQ8U1ZZ^MQ(6)C
PN8%ZXXVQ$K6Z"VG]AJ7 ?7X\Y1[#+*N^7,/27%W.=H[@E_R9MR],]GIMKC])MYEG
P%O.!"[>:2#U?>*8EUD_]0TC)I/PD3RRBQ:X*@Q(113DT0K[7N^!.F.K!4N'//2'O
P:LA")E<[?AZ+JG_ =K9';UH7K.^)! =%L5.T['6QQ<1,NZ<MF%RH&!JM./0HACK)
PGB0:J&_,J!8A!3BKHE@KG@B#1$HG)#E%Z>=LL0V4Q1\H&+Q2)O?[QMQTU+FK<1(Z
PBCM'69!>T'""F]GVC3KZ_X%6HQI6-CHO[6_\M'=OC;&QK%AEW370A;\W2[+S.SJ?
P)(LCAF!1B0C\LH45^)U750O2K'HM8OIN;;W"/P+PY<"L>H5BOT%;%;NGD-D*)L<@
PPYQ#DRVV&79NS&&0AW1_M$VG#3F>,:;E43YLM1=\5T(O0V8&U#A>ZP^9+ELWO08^
PW7,;6.D NL(ZLRCZ)4&^QL:?O;_7J8=F>:R%$MD!;Y@)RSFVP;ZC2CBS[-*BEWO6
P0*+0B[=^E;8$EM8IF?<H[SU9\;=^/,=%;36I!>N^\1Z>*UFIC"H(8DWMA=$KNEW0
PJ5=J^4?*2U#F@74O]J<RE&<G!#-<+B.ZWXZ:><*&[V 7JF'!9>XW5&:8;@,@]G)8
P<(ZOQ?UP?<AFZ)(!=-W2.82X6:I'J=H)A@>!U9Y%(O!(<BU[B^1VOT$A&&FP^G['
P9A6LH !$*DV_![G_ T!=7I=.YDV<J&60Y"DV;SZ^XGA((OIS/G.4F7BFE'2-U!T(
P0_N(5,T^.+WC\L:6/PPU WJY1S;N@COL)UY'4SNFU>QG)%E445>FP"M&)V/V^]SR
P2=X\Z. V0_LM,\>7$"U6BW_[TQ+%P&=@JYTHJ<@QA=N393JJ?_]\G7CNT[Y^RU5#
P0D@Q9GWCGA:^5F ]2C35 B/$?3752SP+X'&GI!O=GSW"K"I\S]I;=5,M G+F_DK;
P$A>MAN;E:=F6X='A\N\<]_'WHA^R]E9G2"]!PLD37'"EX1WC8&H60=X0I58&[3%8
P%*IYG\)6;DHMMH4&\'%9*H9V)?SN. C GQH,"IM:YM9HNZ7<C5I-,:RN*PH^N8G6
P0-.-DACBL\_D/X)_&D-"BUM9 XC"+7,;H'6=? 3Q^2M+'0FY41W$!\B%(+<.24[1
PPKMZIE"C<LS)P@NZM&7A9+XB]056?\E4?BU77,MOAPL5CTH_*KC(B:$*C-ZHF&N5
P"2ZAM8Y-RHI67? ;8P:*%YT3"FX&RJ\(=Y@94?M2)LXQ$9%9W>Z(42@!5>F?^!NN
PXU@%W-..!@EO)0W+L-E]."*#%QY?L'DF&O&?L&G! 4W4G]!2#F\[Q'EW:-3VCZ$:
PBH1TM:[FO3"2681.I$K!R&GCD^$(%/@,^1<B& /M>!NP_3VP;,/=)T(0.8X'YD@G
PT?#S&$;2_95NI^&E-GE/N  N<;,JIX2@>+O',C,VW3X\#"#H"4 1:T!Y46:L3A-\
P.=3%E!3PS3,84SA36-7OP6N!@%\EH]"&;QC"*EH[<'>9",5-GZF,6P.A.K(HX//L
P@6_S0%E\!?+S%\HBBT)6X.F1W;59L&;NQ++"U^J,BIT*?Q38./'[5[NEY2_JIW:6
P=Z!A8G;_4)2$OCQ81>^]\$%Z2'DC7PCB[6FNGK_L6TS#D6I"4ZZ:W:: 7T*_/'N(
P)7G4)%,6Z@N<AS+='67[FK"%RZOBA++F[*].G*U\&_7-6_?<%9;LL[-DX!@/CWDQ
PF8TB,#-R'WB-J62S;KB#()CFRKJXMFU)Z4<UGNX$<H%U-T6>H\2')'/2V$@Z.Y<Q
PEA[PS/;=PIC$<HAV:R#QVS?>FR6B,0"INCR_NGK6$72I-2>-"DP)KL4I^72.Q_/<
P;+.>A$CNX)<S.GVI,D"P+-F@#HIH2#;3 4P"7*'FL#\5.2N%:#2(%3=C)>ESL0QL
PC]19E'4+(5O=?MX>4S/F)HX\U;^;_IT-,PFR,;IMB/ 3OK_YT5U90_)1-' SRH2J
PVI>_W" $7@H\YDUC&N$47 $0H9/6IK+CC9.17$(7KK59QJRFW=]KP>9!;>FT+QXI
P/?Y%L76=FU&A<OCC[;5DP=))XNIS>-(NK@?H%#"C1V]*Q>DP?AHUMF-0H&\1'P5)
P+1!85R*\41JZZXA [(Y.G4PS\U;S-E;./-D4C@IWP6G%];D+BR0O25,9%/S5]U/R
PQ=G%*;C]EG?/$6_><$M8II(JR4B),O4FR*M&NL?E^^K99^%11M,BW=(/!P\=$C,Y
PG9] "E++47<'Z!V OX"2P7WT;-V,H+AB8TMB#U'^8N<TRU3LTMB:Q^D27YN=+-UP
PE_^#+CP]6"U6CTE_& AA5J5T%)Z)[,5FSW#PE2Q?9C/<IOL]GE+CO1\+<'2,B]=T
P@Q]EV6L@T9L2Q-&R;M #O=]KK"+\\YUYP;G+V;CX>LTO@+H-\SC50M8&,F&^@>A>
PPH,K!_#=,U%XG^E2:ZP@98.W.)P6E3C/27K!KB;5S_;/4O#! ]6Q*].^6C 1Q_7_
P47*'?<RSA:I72+Q2^YK-@<VV^U6%QM]*I@+XNTX%X4E$Y:*>8CWO8;CCEJ#8S1(L
P<$D43O< 6UYM62!5B?%R-D2*H)?8JX:OCSMCJ.+QW&AXAX,!ITTQ!8P#[E(]!PE&
PL**KV2G )1O-FW_:"ZZ",\K^\!^?U2&*$W!YF5%>G!)IBEN>T>G(IF/ 7<9VB4T@
P] R9'KUF*Y8;V2(C2'30\)#2D81@PAB7/XQ0C^NO0A+P08"" (F&/OMK!YXM5YN!
P&4^N'"V3S\$,F4:^\2=@[M$V-[3X9WTW%VE0)J9V#BY2]=ZO(P]MTH=$E;VZWS5O
P:UC%I8*%8/)LA/7UPO-BTM3ID40S\ /N"5(ZJKS./(#7EBAACYKH]S^5X@>IW4(1
P4O,'"&WHV'S[IU17H9?+S@XBK-8-PL2FE]RH*4 %!,J,F60N?OB<M/=N42DK*=0P
P+Q'\79 H%S07>_I!MA(RH[C6Q)8_#24Y7N;C4,O6^&?;9E#5R*76] U:U%PD["IF
P%;15!O/R 4B\(CN\SPV@-&WDY9O>;<0L:HB2ME@U+VDBT5#5[_.[HDS_213N^;:-
PG>V^KH,GAJ2H,=4NZW(1X?SH?K^9F6+G,=$VT?EW3_E_BK$!#S7TJE?X:IZ(]A$!
P1/-?_LS@N<.23H[E#2;H3@_T$)795E8209V;#N K2"2$&=YU/!$N# HVD39&*&L?
P'C\7@H"*V";X5Q.H=U,7:XBDR=?Y&C.XN18_OYK"TUJ=O\ O4?Q<5.#NJ78%)=Z<
PR"\WMPL7U8.0(48E5"^C1F]P[5',+R@5^F_OO]8P4XL'I.&X'-YCH_06-BKDR)NO
P.PH5F(3:.3PC$W<9128R^TF;#1T9@=Q&9ICAR9G %U?'14@^%SLA0():*Q50D$*3
PZJ'[H*)?:ME/,)JPC= H,@:S/@,+T#4F6:@'YD2D][BJG=@E4G,DJ%_]+[07_8FK
P.ACLB%9 JE2+07$T'*(6D%*\37[ 4@157V_+@-Q)45TAKYH#CF7LQ$<"V@7JN?P:
P9FLL;=)>_>6M."(#4[F1M1Y,$A"2*V(JGY4CP>SOR[MJFW9/D+_<RS4&%GCY1=]R
PI)!AU<3LP$SS6NE:"EOK4)*.#"(KF@[[VR3DI-!/;1-ZBJAKVFR#O*^=-_=5EU<:
PH8 @SD>K* ,@L9NC(&'Z$'-*1/%V1& -(;$3U=[AE']*E6E"=[7HHIT74+8Q7K;Z
P8+\IO_9]<U6]O=<:ZM]E.CZI%?Z/H[<H=_-8Y)"1_Y[ '->W7PY&\(IZI5S]"X3@
P_QP^B^*):1<7$+^7GP1_+:DDM "0_>_69!7;9JY! "_]&')[>ZP13O[8R&\=5@SJ
PX\;]+@57*W5")XT4/\O_+>,A&*1]\,1);CY+=L1VN;/DJD]O,"Z2(:M_(P._%<\?
P/TC=#5FK@S$QT2_>+(RF/JASB^^_0W>>W$5RX.B)@B\"XH,V$[[^QJ:H@$9._LJE
PX%EX5F4+,"9^ZX)K]2?8,YCJ8WE'R.<"DGG!WM;*%#;*8YO6Y)PR7XSDN28Q"YUB
P_YH\DA<4'+1[LV- <(7Y&T@A&R)>TMLGYF?>BANDCW/VHZIBC[V531>J_*<')EP,
PT^K4>^G I>7/!WE*B!:J^*H1"@XQU WXY.NQ%C=IHO6>' 2Q OOII+Y&%^T8'/V<
P&+GN3!H$)59M/=!*,<4\7P[T;XX0+?W:QIUCWLFL<-N96)&"<Q$=LMAO(Y=-CUY4
P6$OB)R3B_%ED]1CL.:T5)L4ETR/KV\;61M4"3OM"M1[_IFSO'W6TS. Y\V<NS5N-
P-$&?.3M\NTGQO#04/AA#(>S39E+AH_TRCH'M9GI,VL!!]><]'!.#%LEC1<L-,N-G
PL'M/#/R=2M2]N 5E3CH*-+)G')=5^<HTG[>E2?ID\.O=._CDFNY#4&U.)-]6[[VJ
PU.JO_;->XD"Y.MDZ"2CV# ]]&*F>BR,4KK(#V[N?%GM-(:QVUKN01J29QJS:AN*8
P1%UNH4W/PY2(WCH1$A\!>"=H8C=$GF$_(Z^]XY@^'$"-K3<=F]'+("ND;DK.F1#&
PV(ZX>\0=C;AMGRA?<E5ESVAZKZC1:1B< 7*U4] 6JB22L 7I4;9X^<(Q!G592IUO
PI%ID$Y&OZ_.F,AJ@!4:!IQ;RK=OPMFU6&X?/)E>]!%.9..:&Y#G&7PYI$O=>30,"
P(-;*'/**R%=:=IODR_C9Z^YQVR8Z!QX;GL9[SP/TF=AN&G@C0=^Y;M8$_G"EX;1?
PZ/PM*7$8N?;TU1G9^U^U%7#9^("O6_T8;5SODV\0Z0 OF&R\T<ED=N3.LT0R_AT6
P[V'MQ-3E28..-65W:#7;%@[T=/&?476[%'6QIC\38=&N"5U&BP_.F]02]X2:3IH*
P%QRU066L25O\UM-ER50QN9=;\P;C#6&LK6JL\@M$=0[XP->;)_($(;89OV<PW5L"
PAA(/IJ5)X5F=3QT8*W=/Q'.04%IBMR02SN1@D+]$)^:*D#Y_^Y\B!)Y$VAWLVL.=
P!\<$_V'&'LFA%/Y5C6M"#8P\!,?"HBH%;HV&6ZA/;' EY4T>%EAA^)-J%J4-CN5L
P/=2'*BHR0WKE<2V;@!HJ*Z^,IF8 &/79+,TH3B.!GU%E.T9**.PP#>G#H.?Q=_-V
PJ%X-G YMF;_8:C)'NN9LA+/8R*$D#HR[<*:ENX\4'QH39WYCW*5@'A";647V8);'
P(MU26O?L%YUB&;5W,H^[SX>OB\39&;;\G,'=1^+>ZBPE@K8Q#VHY'K1 @Q3HW.^C
`endprotected128

