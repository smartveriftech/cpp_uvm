// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
P7G_;/CPW\,Z()ZG<=X;4 E@3@A&5@[94F4)![=2OXE8_CBM2:R5&$32278 ]D4KL
PR;TFMS"$4GY?M+RS1@MS8WS4'E_%HA &8$$<"2\7\^,'[/&KZZ<S4)H@=@7K"+*]
P^5 &%5VU4V:$^:](U:W B)='N2H(5;D=0MQ8LR>PE M%QVVQ'\6IKP95)T*$KTRL
PNP^.L8FM)G?LO%4T^MN(&7L,Z@;[2_XB7%;*Q@(@KZE=F?LSY$U0YA\3@L!KF*"S
P5R4%^/,/P^0SZ?8P?0PO1Y@G_/!;:\OT6_E?5*[.DT2\Z 0;S@I&DUH]A(^!&Y;2
PU,;E]IMU@_.T]!0;1;^WLK2>SK8M\5)'/W9'Y0D04I&(PQ.2-4C:DZO)E,'G,.^J
P60R/25)5LDB%.-;&R=J2],F6_,3H5F A)FC<+I@A(RH:N-_5!LBCK]FVPQK25_$1
PICN'@TG,L&X\MP%NQD%EEM!7C_QS,?LO-N4R&/T*1;QK(.18O<F3FCM ODUFA== 
PA=N_SG!MJ@[N-V( *W[_%PI3H80@V4)*S#( 6IO:E5TAX>QG92!SBF#^VFN5/4Y%
PS8S .=4Q1/I$APA<E#M:O^QP%<SW&UC^UH'Y3DX4/O>61B<E3X_BQZ!T)"HZ/S(3
PP][.X*1H]TX&0IQM<B66&V>C<FXB-DHM-1R)=TL$CQN2OT\^M6ER//Y=6:TLSJDH
PNVI\U\!VE%='K!H.LDH\]ON""^:UY@5DI!OC&<!MMY#'1YH)',.66I\A;D='ZZ&"
P('T'4S65K)E<O>?C^^P[NJR0',OK: $?&-T/@5K@Z+_5XKE4BS.= 5QI^8?4:7WR
PV0]W!@W9)>.$,:X:.CK_(?\D\06TCW(QU5*0Z5-Z'1JZ/K&W<!WG8/)/' )^WVE\
P.V;]RZ?G[9&OM,WY4R1*RI%NQQ/1HX@D),^+@+VPC4[ +GCNIQV9)R8L5W.RD(:F
PDW[RWRD7U]'V(F:XAUAS 2>OE3]A)I 4/$,^- PK>U/Y-%F*$9(.BDR3F\K\I-DT
PEX"KBTGD'*NN8%Q, W5IK#ZLO\;7(F!;N:?&J>=R V>,"R^V#E?GW!T5@,?7B.S]
P(N\1"^V8(4Y,1=A2B^^]0V&R%S W(8>*BF>$Z6/8CG34,EU&?,LG4;VF-:[C\MAU
P <BQ 5%?5%UWD?$_X.0K<])J*L46(62UF(4V%98<PMS<KM'TV44]&JTFV75\1D":
P'F'NBN)>HI;8!86;.F2%[=&RELX33)>JVL+9X?>Q^;F].4E3)H58]O!A#:0',60[
P"4C&K8I0-G%RL=7__Q6'BHW23W)J ]Q]D2ABEX9EY* D9((C09;5I!LIA.=$'=%1
P0\!":V8UQO9:"7/'&Y*% 6T@*))@F C3UJN!BB1ZXR:@2,:#X_*B6S>C5E[A9_PG
POM,Q])Q"C!W*YDU%13OXN$+-/H"&8;0Y*[P[%K9&[+%ZHOQ#/06UJ0B($%(B$'SC
P\%K[M_[<:-E_R"/]1B!QK(PY_F7<*!*AR&_U8P"0EYRUGH'5,&50^;@=L+K1<K96
P+  #2TMI8&@$2L^"1; G&+MD25%AHV%(8/NO**(Z[%06?>9^$N3>10$WB)>10*Y:
P77<H"O<BI(Y]FL4/ 8?LG6I:T:,"V>'=[F\4/@!>%3H%^HTLPN:3"HAR_7E1\A/Z
PG2O\#7<'=WISHZFQ6M;MSCVB2.EA.-,N:A@J=(/P(S@)89DA1DC_*GM]O5(?V_-$
P[9.D_Y(W9 HK#@!23B2BO$H(4#)KN%,A.\^)A9$).1Z=PV1J_]L$!^G!R9,:39F6
PV7 ^B]BF(A$W?2?Y#,LD%CN0FY7^%=6#B!_UPB@6&=*PU1,+SS'*973-Z;J7[X(-
P8Q76]0!,/$4Y87P+E9!79S(QVLHK("C0&.09').ZJ;\TM*8;;E%]?TC/OQ <EYA4
P&A__%!UQU0:01"FMJID)\\\@F1E?!:=OHZFH""= ^RLFU/7M?X C544Y)F3%&$ (
P;"19\,04F'%7R<.,5#3\E .DK =YBF%X<%FJ#+XU,)8\;Z5T1[K]B7H"8&MO^U%Y
P=5^K.<K?#T%BPW8-*2!@\L\-1B#24;V%C2HE0W@CHY04>W")+A"',9=XV7T%%S1M
PH6!UAO7-PG7<"M?):LX9^7VJ\(-RX%3F+? 9T3(P*B[6>'ZLR-)Y:O^%>Z/UYHB$
P5L>F'N<8Z2/@2W8N7<UN46T^Q$FL9_7MH*FQGM&JL8F01M$X4DP;E&'@<M05C%=%
P?9+^$;$D/KWXBE!YFIDB<Y73F,_:\LSS<2T2(Q;Y"H66M"!+<U-/!SXOV! ,Z!VS
PJO%#(9=R\2K<A(0[DK*% @_B*3N^NGAO\2X3E="QC>?+%/>:5JR\- ]A_S2J2#BG
PJJDXUS Z4,BG:YRH*^-LBY@+3T"B;TN!?LWZK^8"LQ1[&[,/%<T,8SW\X?^I3(#P
P99W*$A)^@)BRK6E_'J-Y<3+,/Q,BIG6=*IQIC?O_Q-OF35MI=N "!#96\818NC\5
P R]$?)R7XT2W"NJ/*D*SZVQ&T1ZZ8C0(G#35 VX0..\YZ*YZ#A-83E_W)$D<<0A?
PJZ):L3=\E,S;I45ZYJHC6 P&6:IBG028DI4[O*KO4S1"XO(+THJ82OU.9OT,E[PZ
PP:P3UMS1NA/+C#1](0K+ZY)[1^/L*,ZA0ONH&\+^&<,CL.!@>A3[/D,OGSVFI%?#
P)3BP,;V/Z9F=)*Z@JHEYGC@(HE E&3MCU[(K>$BNQ.!'T?R1\L2-5@<21$UP4CCO
PR;+\/5J/H_Q[[G#U?UO)&)#:5&!Y[\0R_P"@V^!JEK0N610HX2/6"E/"Y*](&1$^
P4 ?4.7;T#T!+!:@9T7A$.T<5B35?T6%<?#U)*OD?@\.5"@H!7ONIML#D5[W<**Q\
P:5*(DOBN"^(K@2\B[@:PTM&U.PGO8'*I("46/[K+L(]IETL"+<'O/?"RUQ#D[9<?
P2VIO; 7B.>ROX9>2'L08N4X0+)Q&O9][EEE721XSYU79<47]0_=_8&ZR=L"<F_"!
PE/-6'RHY[B'0>CQ^4/(?K >[4%3GD"UU?J1P.05I<BG$(_S63Y\=N#GVRJ/O9U&H
P(V08K(?#U]K38G2Y(<+.XIW>T9HQOA+ZVW2DC"^K. ]W\@ZS]RV1C[EJ8\755'"]
P%2/;Q[M<CP:A[KXE\Y8:@95E[;MXHLPS/7'=X=ZN*! HKAS('UR62SWC]6THIBMW
P?G$9SSG(VQA:9JM?#R^H37%)'WL1*SV+*_&)@1P!?N23;&]C%!2C<<1MF*IA2;]\
PMJ9.]:/+%B)/]^K.#399L3;L XE$^M$?^TJAWXL*[LJ"N4>>B%TD5ODF6PY7'_5/
PG7A_J#M;="688T 5CU:L#:%.CDN+MHZ8=.J-3^AJQ?VC#G_-MDD> A?3]H$]KM[$
PVDW/!4"EA RV$;X:]*#)S1W"9)N#?]-<]$(@ 0@<MS+94( H((/KIZR'<$#ND.;:
PH(',U*;8IU'Y(R TGH^4-9O(B4IX"#F7VRFWB;>>2WM^UG'!G'^-Z:<)4F>9>GT#
P7^:!"C*N%K.T0QT0\=*[!!J%L$_? *! )D*9 82[4@.F)I5*F5-NA%CD @%WAU1L
P>/5:EF7*V0)3ZV$MV< E>N_32;?IF%HX4)58:U=8QY]Q._?H$RVMU%NR16A>-];8
P]DUR13A%6O,T8?>Z843KV+A6NC,WD#/+ID:2E_2L<IYFS7NN2Q.9+"F^OSF#OG;I
P-')\:S6&*O%:J'6<,)91F0EZ]+G.*)MJOWI#@_]6@@2M5QV<$IO="MB546E+;"-&
P=Y7^'^-YA,>&_7P!4ZLG+2]MC1/],U7^@A_$7SNGJ&][ZX=CD!_[:,/ZU7-K)5.A
P\02%C@E2%Y[@BI4VJ!T8G1C4TQ.@K_Y58#@YZ5?OK[):NQ;ZV(LY-Z5?Q0M56$^T
PS:R_Y?&NZV>*)K\<1/+0B4S!,PQTN>S(X[M$HD/R\^ 23!HAUTA223 V)U 85JE+
P^+<&Z)=+[^>TAHR8G,T$DV:[]M]]?T6+#VLCB.?X1,&!7>I+Y4_T61>R=#"YW&N9
P1':_XH:;)AI$4:+T?S4\@H'D;<'<2U-%3MT?+RNF%UB@"8(P_,\B?N!R#<WO& X9
PO9BYP[-/<'O)-CU1ZS(![-@EG0*6HA69&A-G5OHJ"$A*>P7I?MVTER/TH\&M-?7/
P*LJU906"C4E-ONUG:B]5"<9]EC<0+9)PV%5F:$1=RG^?&(5!(#*'[E>[G9N-$9NH
P-O%S=1\>SMH%J\+T"?XZ>@QGN(8W01SAS#M68[WO_>B>9C)3WBU0#?$-L]]0=F9$
PLX/%6U9=F_397P%N5&?&E.R^&W#Q\C# 59.9<\7A6:-_X)K@:=^E!LU9C]2K5LX.
P;'1]T\'*;[N!%HT1.V+'!<5JX2M3.42SF_.CRHLMBL&'9)L=NI5$/RCMKXP>VVG8
P!;6MOOTXHQ)Z ?I*=6%J/445/T$0KGY^/  9JI+AOE;!QIBVQF2VPR2Z[L:2J>##
PJ(DO,>Q72*ONX(6I:FX=>J%2?PXUX0>25Y;&_/Y#T+&X6A>:(.&GO^ Y<;G/(4YH
P#NH8N P4RX7KEY26<;CU^Q8Q?[%^LY$PE<_CD Y7YT[ L=<2,C[.:E8ONT8NT-"H
P/GG7X]B>?L9M$KY6MVHO>K+?,"FAQDZP]3B=> 5QYT0_@IJH-U$MAPSWTQ@+V-"]
P=#Y-G[4KB#=!>*8//'\,9T@OWN7^*\I%Z8=L\KY%Q?4:MYUK'P3&QN1 %X*HU(0.
PQ',V*C*^J%:S4&C[6A:X:*"61ZL)H=RI*W$;<-DCSQ]<TT6<W"L\=2%SQ*KR5&5 
P&V/5CD>EK?@5OJ$Y&VDI!0R>\"H:R!)#'<V%IL)D,Q]G25C)>#79%S?G&'(E"B/"
PDNQ9,#BV1(B*D.;#94%Y9 ZL0@_">G=X-3 ']GXUE\E<)'OVX"*26*%<4Q=JPXCH
P$*+5CG$E3:OQ+W ZE3<%9J[:Z21PC$ M_IZI8R;Y> <%^+F.OR2:8<U<<+<(@^W(
PM72'3^FJ!B[Z=F%]SODE8(4S/%UPCW?*%EM,:FF^=!49HVD*L-)FN?,@#^G;W$EQ
`endprotected128

