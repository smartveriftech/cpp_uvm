// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// File: uvm_dpi_helper_base.svh

`protected128
PW/U^L57$QZ7NA0%,V"^+=&47]V^)1^ICP,/!"4/LY;I)E-0C--2C^#H=OSO='8UZ
P[#B%'./ XSY+8'G"W\PD:B?&_',26W=\*"H/\DZS[\$WQ:7Z&FHB1=3BVP/G,^^/
P.,PPF_#V_?@UN*Z[,B$@\7Y7L\8PI>.D5JB'5:I"D9%FDL1AAG#F7EEZ0;#[7U.4
PW[15CA:'*V5$1J%5_S  G3AJ\LA (3"#;Q[LB_:+/ $!.Z7^FB\G7%'=9\!(0?TO
PC> #E>O?9]N83C45>R-R?@HY8D1.%^OR#3]D"#1<O8/IE'@H&T]Y>0Q9+1FVP!2$
P7&:'Q9!+'H3Q*1_Q4<$$S$??*E0?M^'2*TJAR:CI'OP_'-3X+#^9/**1ZW DG4>T
PP)B1MFX&%II+=)F(C3$$H(+L*R=.TSD')]VU<6ZA31#.$]DP-J@Y\MAQ6]N&^JQ'
PES44"Q>HZ#_@T\DDW">+HFKAAC?&-75D>*^';[,1'VLTY/E:X&*91D("[BE*&_1Z
PXG^K6)>1!*PQ""?RP.%O8-QU0V:\'9^C-63[>-SHS_#.7M;>Q(%T9M>%ZU'<LH],
P-KO 8?=AA._&)!7%3 #HP*V8312)0Z3$P^M'91B8?]=Z<D0?7?R.G4N?*\;-)W]2
P3&?537:I2$4R4E?5??W83AJ9Q'_O@1)H1$C&DQ5*)0&2Q"/!/ (SDYW(=S#<FF+K
PBHGO%BSZ?JF=\)1);1MIAQ62BA&Z 3((/&PT-0Y=CRF8Z^@EF0_2E7HC%Y:O2[IR
P<FC?=FY/&GRUK%AIXN,J.5; 6X/WTT#%9CUER7[\/?H14[4VLWW8&*UV,7=34(OO
P9&7Y*45\R67A_#03P=?!QC578V(_J8=[?FE-2 /B&@VA K2%C:YV<2R^6.-$&T+J
PR0J"-(JM>705'2T('I4$5W^0F?W90'-I;@<'F1E;_QZ&C=V0@(FLBH);YW%R(4+#
P4X@DQZNU#XJ&=<.CJ;VUT/(GM7K'=LP]3=)I2T>Y^5S!]/'>NS/;R\T%19?6,!7M
P5-9K40%XCB*2($EBI9&\Z_;%A7@<*SH)VX];-!A)H*_6]Q<<0#G6MM0[UU1:=5\U
PT2K#FX/MT>V"B53DJ\G\6C"8M> 3[#FK1.)X962C3$V1M$5CO57<V1)A@@X?[#<'
PY!"B5^@+!L'\$"/>P9Y:736ON#^']L &*,*;-L8SSIH+#T&XBVSE*8Q^/S*WP4^L
PM_.""[:S"&!R5"QE9?556R\2QR8F(5'W^^!$DV,39,U*T!YLIQTHXC=>-)V9^*D0
PE7OT(R0E*I=:4 FD0Q\]^1J<!J'(BNN^<6QJ#:G264=FZ$WN9BIK@="58:2EH^/@
PVVDJ6:,E\3  2#DA[()2TW^WB=[\>-5&<\9D['FB&O%TST_AM-]E7*I/U>7$YWX^
PY%OA\6(=S#$\[;-@D5UMS"5H2MS=%Z)BSXE5AD5_,F U4.G17FI_C _Z[+!M<\$5
P%Y4/P5=9R#3XZ]F,]LO@4.?]FA^6)?>IH13$63YHV#]$[W'B$;G-*7+@LQ^E4^.I
P)A%TA&5:Z]49D'S85[>R 0>J$9["C+]OW*Y1DF?9^:-HS,<9P?]SDD#^S6(C7%CP
P$G_;%.&F\6'\$A$W.(!8*X#P57V!IA?TH_'H2!V/DC1[XEJE<>G<[D3%?5]-$#8U
P,DNH8SGQ#KI1]$4^=#$V$0MJZNI,MT$%PKMG*6+?<9;2WQ0'&>S#,FSWKU;*ZFZ3
PCP$!\FNQ0\D;1U,14VXT;'7N0\$8?/!\"$PZ2J1"N*'9_]! !A<$1F65*E%GS2)6
P_F<%BX0%#$F"(_Q!,@<*PUYW;)90&Y^:ZOA6S=?I5 &R<7HLU/?QOR3!!DUZOK+/
P)LY.#WI7=.I<^W[R6>8O/J7[87V%S'/GHCT@+>QF[*1;75V)N1O6I F$LIZJIBH:
PY(5[I9RB]-5FB::6^R"$P8"9Y'L8-5]-B>:CSU89K@OBL3$V[^7]=. &1J=Y+H;Z
PIGF^;(7%)=7A +U6QH5M%[MM*V5%-A<O5DM9TEM'5-)XS-S1BYS=J]D9CF7%"5*!
P\BV(1;::\C/6-I0N'LM*!9?('[.H'['@:^JG#H3%$L.Q_^T3)MNN].71M\Z#XR2!
P8@+%)U_T"0(H1CIMSIF\W@O1FA;E+C)0&#.3,CFPSK(ZH4RK+W-]HJAX,!7;!I"0
P<T@.&\XJ>H'T2NX(JNB6&,[XRT'LGS9P#\I:5CI#72!V:&]DNHSU$IZ1L!W(6SI5
P# EG6\L6!< [I!$+B,,U51UW.5IT%H\)EG9D-\N#CU803[<!BF?6R\,ZH+!7*DNL
P#_H2:$B[5DJ.H'][D^+IKHN^FV6!"BS'.JU*V; ^T5%2FUPP(J)-'YSDQN9#M8H;
P4)'0>5N<(J&Q/K63V ;RM+0"1QX#ON%G!6HIA4ZLYLC^9! +4#XJ!ASR)7 ][$-J
P4D]MM>$"RDT4</D-&)- [BI39)B3:>7?(YI%26KG/\&Y*)BCCB-$D_S4HHXZ2>6.
P32<;H:**WCGH8&$')=P%1/QB^!*_(7N/WI_NH[*-5]=BJ/\B<?-R%1Y[PB4 BYQ"
PR%="UQ'D-RUGV%-;!;Z1O-XGC65UL6$9?!S&G,$=VM*D,BR-&-J5JLHCUQK=' M5
P2,B9\'6PW;<SZFV?HB%RLJ<O&MN5;3K9Y#^DI&0#$LM X/#M4_[+SJ$=M'P'#_"(
P4XTJRA8\.&"_]9>LZ2<(,3WE)Q:_:+H-D)OA9P$[_Z7J/J:TAOK;3S/C#%6*K5QP
PK[R94$/(?=&E>?4T%<HZF5QO[I6USYF$<E@#A.!).D<Q>"TZ+ZU#GL.P^#YAQX=<
P"(P.K>L$3X'RK=&FK=KC^ =%.,">'C0QC#-E2@H$T'*W^BDU0Q%ARR65#Y80T7 J
P(U'$;RJV:!$8D^K(M3 F4AW,-*N4!0Z-[_V5M/6LQGT$^\"6QM1=@Q2 %>/LTG_B
P0,1?V.-8;,B]P!4.&A-^3O 7N\*@\O_2:9S1Q&B30,FF0G!$.K97YD9"P54_UM#?
PLU^['+8HK[10VAKALA,B(A1)*I0)8(UF$_!C@+81 ?@-KA/<1CR[2Y ' $L7T51H
P8K?S02^#QO!?L%2I>BY?4ZYTHXW9M^#]1IWR^8ZMA2N0G%VGR5\SCS@VBKT#FH4A
P!'SREHUE;\G"]D!4K0Z<?8<T'!:HW%=4"*2U(=1-B^*M 7+"QDH8[F"[G+(<O"6I
PNETC9$;G!" 7P#+MVAXO&["U[D99(WKA'R_D/V4@3N[M&)4,T?Y%TS(U2&B9!O^:
P^N_544,$ ,+T7TA+8JP@?()CI,M3 E79\FJ(:J4Y_0S5MK.T-NEE[P,YS$Y.UK:I
P$8B?#NL/G+OL!(-/XY2X)BWL7E23)5:QK:RH?2)E<E<3YV*VI7F;@](2S!&6P0R)
P)W,/YH^9%]NG\N0^3C-:X GB(!NS+0%IT<G\6^!6PH"0=@UM_!K]^\(0U[L?W2U_
P#N>V#>_3#=7H1>9'KQJB'=;P%E%06Q\$ZU_-U5  G<[?OCF7KBQ$2QXYHD>WKOI$
P#?:*;T;DRWL)POH<%2UY)<TT<U"R.XL>U1=FF]#=+6.H$AJ67A[D1P:E\6#V:,W)
P?E3*G'6"^6M28/U[O:@,]ICCJIX8N*.2Z.'@XF_#.2HGF\Y# CQ88I0KW#>0!8*L
P1.K*4'J;"2Z'?!V+AZV#N _F%^Z&,LJ\@J8>)5.R)R/G%#O'X',+KP<6/5!7AVM+
P\Z;UH44UD</_CN%L&8JHW#1/,^[67!&?%=K/(-:N)GW#+4U$PH*_2'//QEF+4)O_
PSM0#Z2;XD1'<.H%%$CB(8A^/M0LLC9(JXYB2$L3Q@Y!H@NINKS=+ S%BF0R.6L8R
PE.X!5!-BL0ZRC?2I:S(;OCP6\4EBJL78AGU7W%3L<GJ%2L-%7\LU3N>2_!VE(AM3
PO.Q[8.+<?Y!RGNJE/=,8RE(N[K8)G":^IKXI0IP*I(5&0X4=7CVTNT6V@FNE"&MD
P8+@%>&!,)4 G]N]]+C1XIMKQ"F1N(#]503(7)RDI<" !5&QW*5:P,>GL]Y21A?^Q
PQ9?,UJ]D_TK/V#$)J5VO2V0_&XPE /^QH[*L."(,M_>N_&2B9' BIS<%D5T&L;&/
PSX"_,/,\CM-&B]YW9$:Q0 )$P+IS&/: <H@-4(KH1(*D4Y#D-J1@+H1^_!)>:!#'
PTUU'/MH?%-CZ$!B6O@RWEX2BRZ&!63:5?+R8!S+2^P-M^"[&>$SU*!JCB0B=2LAB
P^#G_(EHS8$N'P3"99RVN+SL_',6-A1D>&X =)GB34HM6:X'*7_WJ3BH;OFM? 'J$
PDM1(X8"FVNRLH&1FBP8O-$%Q6UL]\ Z1TL<N8VO'>98?12YP& 'V,#2D95J*%%0M
P;T>#T-?LZ,:6XZ6\7IL*$3%N\7BCC=:[P/4@="<-W,3T_I!?6J!CVQ,I#&P&PP1I
PQ.0)-6-U+ZK"?"0W=[$>]!132 F9TG!!CMI-6O@.>0(UH2:0D!G'%W4=>DH0'"(M
PZ<HYL^=*L52'$R4><AB:]Y[$ZA$9Z3U!DE,WU4_@^^*$8U"1^X3KLK_QVI##[#ZH
PSIG6QC:0><!O]RE&7:K#_^.KL(<-Y_%%O=#Q)IM:DNNR_M:+2[V\NCQ5T2C7Q86"
PHWOGKJ5OSSI8($0FFMX9_V*<CCW.UX,9.L1!M==*CR]DO&H*@\NB=A>[>O.157 B
P#!EHU"/IB7]8DJ]#$NFI;5MBK3'*C1\15AG03AN]*./>!S]Y%&!&/9/"(CJYWX#9
P: "%5T3SM<2Q =&8PV(!ZY)&W(I?]>VM9P*K#/R!"SA,*O-6A$E$> Q5FN3]Z*@+
P#0E)39@+ES>'V3YXOIHV*ZB]8T[2$?NS+:F&/Y4&H(O3,Y#!7G,AM,QKZ3@_0T$]
P0EE96G9JIY_46MD_PG$'(/^CLP([,QA9TR-F\?\;*KMHXOK+$#=]2%::D*8JUEJR
PKB!*,!JB._GG7.()K=#LLA-E@7TQD8["!M6,$'??:QA'**-_2-[!Q>@^S]5LZ/AS
P<J:61=SU211S$V78;>$>^GPX:?F)\FNG$A4,\S!#EIFPBO[MBT4R6^692W$S\>(<
P:%(T6[=50L4B.MK2)IT)5:&*^$L5'3CTF5.02;,)[Q(H%R,'Y$^]=\YCR# "^V5C
PZE]>S_+]XM.\J^E0]?] [O:H- RP,NL"<N23?@8>2P1J>]/%Y[ 6D+)VX(RG6NYY
P*.2OY\: V3@AO!_4Y)3.$H%,N7(B0NPK@!]2SHV\\C!R9IXNJ1W^N_ACQSMHSU/-
P%^ YJ) M2[)<N2]6-KUJ-!*T\+^+TF,._>8% 75*B2A0649H4D+?=QX$,$*;<%CZ
P&-WT#UST9]QV,%W='ZVSVP'.&8Y>_HV#4(!FQ4#0\DWVR+0Z*0D2^3M=)^K2  >M
P[D"GJ'UUAOB/+./'.X1>W]W=VOPE=?$ Z/#+C[?\(TY[9M&X+NXR?L$S$<K815\U
P('?QZK0>@.^UA%8W*]E$E8[P<$OQVR0P,9<,>[0^3:3NDV1A#7 8+P5,QV,I]@I5
P*<?YGM)'OZCV5!S@F_]0!C%X]87O,0E=KW6YY)*5X9=G(R) GV"%;@FX<NJP4,Q)
P,TV&O6 ^MR<L(G>/0N3HE&1Q'MP]5UCH<Z@Z!TF0B K@>ITL@1#:J'67V#/:F=$:
P)KAK2YPQHROQ-91#KG]+:1SE(S3QWZ/)X#FCO\ZYF NU6@H=_"Y36+)5QGVZ03U,
P,5;@2D[J47())@:%[X2\O/,CSGI#&VM3\1*SA)L'N'_TKK096LKN8"E$.ZO='38J
PU[H$]VF+-#=-P[:;BC<E]9!)Y.7?YTLQMIJ%O:6&:EU55856T,8"7&:5_[[BS84(
P)O#7D$+@L[+3Z 2P(P->LJCTWE/GBU8A<\][#)HU?BRX@2<L5.Y/JXYHX]Q^*F*/
PHH;9S?>3ZX0NX_R_,U4T@SFS,?08VB$!FP*@9IOX\=U8AD;A$0GDX1W*A&SPRW\;
P+JC$:C2VAZ0.O: M05L.43^*=2NQGB$76?3DK$CG875IGE#Z,!4;Y'9$9H<RJ85B
P=$M0@;/\PX3-ZC= ^0$B>&._YWAVV9GD)9\C''28#8:E_!$Q"IPG5HW+M#O:#-#1
PL3_3*DPW$59S"T\_4VEV))CGK_%7::J^%''O92:].S*G 6P[IEZ!7W_8JSS,LQX-
P]F:29DAZEJC#B(,^]<X-#SK44'TIHRR V_''4.*5;:%(KY!3ZG11)@^;/S>153:^
P4WD,7$=.CP6OP1W.AV7>'7X:__8NN,M\F9#F.@%C_>JX_+@"247@^_[>J\"P$QD"
P3*JF;8]XWD$=!>Y-T*?M!U*I8V=L6H0.57$@X_@+/#=>7NSY^*^V=DR!((RVH=VA
P*WW*;1]JBPWS_Z'9_7GB@JLD$-^J!5VM+EGG5V=MG,G(]E?6((*U@JY"U_-Z[[_/
P!VRH\K6U-P#Q3T)*98HN^MP$Z0]#W@B/8:#L42H>:RHOL76=?LUN/"&D,.%I3F-2
P6ZFH(&+G/32Q<.?N^F WGNJE'???J<]8'.N;G0NJV'1$S?[WERN)WZ%\R.@:;=#$
P[N2NS4F\"&FC*SMMG7CIC,_!7> #TU+&T++,$->&)'X-[36K=V&\DDMVP;;K!F_D
P#E\(44;<A; >>VIP-ZS=V'6_P4LEI*O2K%1:!ECM=2H".]H KX,>-7Y2>H04.$='
PM+GF2IF\I7/AF4!CQ3;#FJ-VCHPF*Q+@+0F^%8!?YKDR+0LVODY22G,;>F96^#8(
PJPO@SWRY.*,&U3(O15.FM9D?E<J>Q^) D=A,J_>RSN?V8VGU!6@)7._?;3_;*'J-
P,SC[<X1NR1A]B&*SS+2&;_52;]VG".3YIN,UI)QV5VQ4]_21HB%&-FE!QN/\ZAM^
P1^Y"RV>?SQ?PJI.;&8#M3V=H;NK))HZXSC<. KPNFB)+DO]",A%)2Z!J")#YN]>M
PC2J/%>$-*+N?!0&B<U(U(!NB''R=8RHPYCQRG>$L\'Z"JX8Z;XU1N-JA&J)5-@5H
P$_(D0D&B3GX^P;E6)R.$LQ E.]@Q6U6X4Q"_:O43FW,\F(&W?>-S/MM-_/*"XJ?)
P>FUIBX 9\=K2&+_/K#%NX!&_Z>D+ /K\6A[B(490"7X: ,&WHF8-Z*+/HF@<A -$
P!-(K4:@8>'.*"1_.RA PL^FE=3\<B51@D7OB8IT#?._IA<D(,Z1B68L/-HW&@PRC
PS[4*@QI8PGS3WMNWF#TL^06"6M>UQC863MN@M[A;J!(3<S#640_KQZ7;#X;ASVAM
P;/5LX^1EO(NV>TIVM$G*E&$4Y9KY_!59M^_:*B^=7A%)6T_60;+IO3>O:H_G:&Y?
PC,2VK?;U]2?<T I5J_G@,^P<0$@LOFNE#]A8C$93JR>*["^#;:&T=*Y+86)?^^&7
P?;AW=<H%+9 [[!-T9/!@KDOTYMQT21S=S5>8AE#?8!<B]-Z,",08 D!.,BB69V\_
PB5@%E/7>*SV_N/],U^@,9FS]/V"*/(T0$LR2Z</L_!@YKB\W-?ANS&<4R9N]7AJ:
PA9F@[ ,U:+99;O_'D:FER"T=@*,<#FBJV;\>J$"I!-TG=GY8KS(#,Z,; KC+C8S'
P!,9HBPT4(+$%G0;X29K5)Z+@::7!/;1[W3\^<KY&F&LL04 K:\&WK.E+7>6TSDA4
P-Y-F?YEC9SHY;&W>Z2T<M,62_)RS1T#*0*..TAIFGI@#- $VRE#9>)]5GK-24K9I
PI5_XGZN/(>[4_U3PW=]ERV<$><4VV]$RKO2#;WWC/',AAP&=2FFCFY3BCRLN(UF/
P .I3YO!(+=1$'KCD[FUXHJRN*;[:7U)35QSP4^3UG:5929T;J7_<+F<L(IP]0>1<
P:>O+Q[7,<0;)[QF335JU]"O'-&TPC,D _/6QBNE%\Y_ <=!\L!@ 4WT]+D\4.9T2
P]:NO?QP81"]OZX7X'7F09ZP>WM="D#)!BSKI2C9-/_'K,9?IX(]HC%6D(,WN6"*.
PLJX"'CY,PS8/YCRNT'%I%.)YD;TB$_KX,L!QYZ,^,.+2+E+KF+M">((2E]Z&FJR!
P'7M+V0\[H_#,N-_H[2UJF_2P>VDXZ93<)IZC>B(.=*Z7$\3-/@ARKFW<'N"<N$#H
P(@PZ4*0!TDV!M>JM4Z<D4C&?"7:JU&U2-=DI;X[),=QJ!+H\[>0W2PFO[">#@L=#
P\/$[S[*6HG F />';9:A+^7??]$OHY6,H,F>$9IA(GSYC%(=S)^=\N&N]G]6G8Q8
PKC:>HT?J&CK&].R:H1LC61(>I5ID;:Q'H<&$X>[5+M?M02A*!4#9=+4"0I'8CF(X
PE/\1(H)7'<<-UD\C4-[<;H$&<PKV"F;@.KF#]RJ03E(":GK@%U)LQM!P(S44Z\R"
P5MB&6Q)QTX.MI$](=&IPQU,#E,U1Y3#0!F2U )SFGFGD&]5MN#M<4O'[E6Y;HJWB
PNK\R7KS$T%L2>I"+ 2:J]V$&,[8AV[;3&<\^?%<P;6^CP^K)*)GX@DI9.ML=,@VC
PDO/J6?GO8VDTO[>UWJUA8,F.]SNV";?/Q9DUF59JT<C-E']P!@T5/*[YJD \MDT8
P72RJ )@^9WVNQW!(:9Z!RU>*AT*D#&5(&]S+-S"@62.NO)7'7/' ^J-[WE/?EEK&
POF.\W,X$0UBRJ=]HI]$?&\$\ U#>3\2"^31[2OF;<OZ *5A&[ +.YC54HX/:7UJ!
PT$:1>2X,,#>7HJ/YU5GF,:&H8A;=MK2,L!'?,5@1^S$) D=TKO@,**N+51ATEHOG
P!!X9477QKA1]PA>@%.^._MWW^!AJ_OZCFD$ QP"'(P1+;<?6'_*O1@F=6\V\DFC!
P0S7-98;2;JTLB8U:6Y*63+/01OL(\UN0$ QQ3R4BNLM#\!\;  ?S>Z91]E*?LSG@
P[@#%EP]!^9DL,Z*\]*$5N@:$BTM!F"[:U#P[)?=DR:\D7MR/$49O</QM6/5!?+/!
P0A8NVEQ&3K#QDY M_ 88ZFQT>#*0,Z)F*"8COR?0"MNQ9SR'#A(U8V^24.M5#>TB
PBO>L8#ZRCIDV3)'XN%609]T#9*R:Y,-MZD 3I57HPS$5@Z3C<^=L%@RYW[/.KSCA
P?;]VDO4:E=V_G%(YHZ6;>)(71XD/AVQTO[.9@-']/3L[HQ%E)P_]0S+!S@+',-%+
P.;BX/*$R:7KM[67[=:\V-7APMT9W!WZ=89VZ/DI(P:\)F<WIN07.Y^];32K1\'O&
P<=0!\,A09C"VK%IK"&=K)A0D49M9L&L&N)'EZPK(H-,NPZ\Z?;QA-VI&T++%A&;A
P$N3"L)]U/\JW#02<<%)CSQX2A3A-HV,]EO""W[\^>"FA77(_,F*4O_5"KTBZS N6
P8<'>[2'6''DX$'F*[A6%*YH7VCQ8.)Y@2J;.K)'8X4\;_G%QU(RRP).S9"B;>I"U
P?Y#=56MNG0^^K2T9I@^VOBT9K;S(3 LVB9&)@O@,Q;F'-;6J@RY.DS]U%A<NI["6
P-P^SDL"]/AEZB@L=S%WA(?V_X/K-"Q;?D([O-XNI"?<&+(9&HEM#&/03UW(\@5I_
P*'4U/$O93[!#Y#43U&EL8'<3T=-9$!L"/5R#9@#GRHWP2BV)"X016&%_MVB"+HQ?
PLQL@)1=T),%?7O?$"SX;@^ P,%' :0,VU,D-\*,WPLM[UM$QNP*S?5-)PW ^H-MJ
P*=O_G+Q5E(BW.)E*VS692;$BW<JKVYX/*[4\"O>5QJ'1R[?,\.8.)M;A;^";RFJ;
P$C?[$_SFQ*4?N6PBA]ZFC@W"&ZSG)D7S-AF=MU>@)*RX1(^'0Y84R(&+%M\9NEDR
PGVB^U@&@/F]=Z'>.=TYH(\@JGV1$"B(J5:^D28?'#W=9QJM,5NOHC=I]O_N<W(>Y
PD2B#]\+*QMO>2M6-$.TNM1F["7:5E#483G"V<[]X*T\0$_^R;YMAPAM^)V&&&D'$
P+,MQ!/,[^31R;J-4@G3=&$\ :H%Q''7I9W9=-%IU<TZ7ALF]T.L63(#=IQ.D#QZ1
PQP'G%WM867I1VQH"9S8+G]S/EYC":+UVUGVX,!%>U)VGR\I3U2'\MQ&:VB],?^0S
PKMG8'\@6E09RFIN?J@A/4.R2!E%8R@6QV(X2E2/^ 32%,W4+%:50DMR&NFOU=.;<
P5CTBH5-OADZ4T V>MCXKK%MRYP#(B+0D^?<]N#H5RB9'Z72 \/CS7P?1H$.)#"Z'
P@)Q?2B0LGZ6A6,PR:ZY"8GM'5L<_-]<:9SLTKQ:+T6)LZ50I^\LJLC7H)M&.5U B
P,FB;E&9]!&ZZC%]>(:#.K6_+.HJPGTOP@(5H^JC;@IXH[>'/Z,CU*V!W?SB!P$CZ
PB1:+N:)\^ECD_Y\J (.K+8^)Z@^1Z'TLR!X8Q(6;IU.$A1T C6E"VA!!Y#KS5K$3
PR1/5U:P0!NSC]\IEO<L7EFOIR'/%(2:T\JJ?0#1 E[P%K;6 -HL:YQ<G;B/?9K88
PQ6\Y4C!F\3*%_4#9)(W,B@]=Q):L)4S1BF/B&>#K1^VR8GS]+;DN\(F#O5RX-[X]
PY@"DWMFHMWY%".S \B2'^ (D-&H\ORGILYQ4?$"(FGQ20"QG16D!?PMB4:Q)O+]7
PH""D:!]H-$'P I.Y%9+^XWN*)$+ ^$9MD(/&<_-\S%L+">4(4N$AE;?2L8R>F$$T
P2963HEEZ.6E5!R/7?&CC[RLTPC-<&""5<PP^F S7.OSH#MBM=G3L!F*AE^25A+5_
P=P)>_#MZN!BOW$"J$'6S-XD1P-NS(H^;.82(*LX +V$=Y^#&]#/MJ:WH#99;E3F"
P^1T$"'Z.JP/Q[)1Q[:721_&."HDG7[(;QP-1^[9<666KW0DW%VIYD==03+^D:HYG
POE.7BPXR5:A$F8[4*&40@0?)1,8"S3(85RG<_'+D$L(6HTHA83]G%K>84S_QJN#5
P6)Z-*"^7DL"\R_I0C5]3IH!4^LKV48+!7P,8P-ASQO&1N\=W(TUNY]LOJB:9(7A[
P<?#Y<$*[$B4<_<!13)U_O$GB&;ZZF<_6P98_5X@P Z,,AJL\0+^:)$0<-V21ZU$7
PP[)R)L&H]W-11L2E!QTIAX55$4W^@*.W+;LY1#&Q4P!IM!.)3 P'R\]FH\H[A PV
P]*AOQ7$J3!W\?.R*^1J4L"?Y_[='9Y)3QY59II]>WBA ;6"6\8EM_WV]C[JAG8#0
P/O'W(S#)TWY&!AU;JIT,$) #4*\RM_S<7?9 $7O7Q/?ES.@TZ88>HL&@)J8>5HH_
P!_Q'-H+(E\G/O#J/BX'G, KITOFR-8&,_5&BWQ,6;F91IQ;84-GY2BKD9+<L;3'5
P9,7 EA$(N/.5)P]@DS]L:*@_ 4T$ XRVXXYMCP+,0UVW]MJ>)I@%Y:S3,MQ1C@G%
P,FG/@I8?OU,#]Y3+FWF]W_4XR4WMMXIG)2\M?-'(?K#5$B.[V')>@GS*ZJ6=-2+=
PZ%'Y[TGF!YKI1"K)TU  L-/)Q,=VM+8#W3[WGLS8D';?B<=XI 6G"Y>I95C='-8A
PD//RQ?H2O3;'K5:WH8=C@8CN%A1PT2I74MR,J] [I70,OF9]8TH(UMY_,&H<AKN\
P;.M,!SDM7X:M>WMJ94,R0B$ BKJLSP">28I\8^!^Y+REO.^A\J0P^/O2B=M'' T*
P1#+/0+TX1M)Q8,BNRJZ%Q]J3!/C&JR0B[&@UU HI,5';_GT,4U?AA@'C*WA/%%QO
PG+^';,"N!2!B-D'&8U . 'ACN+S-&+J9LA\7J=W#U<.C'G R7NO5+J0D<CR8MN1Q
P<0A5+X5AO]Q 8#YJ!D[,=&N$K)Z$,4<YO/MSP"W"(E'GGU^R0%M0Q.U_@<XVF3")
PA0F#?NVN"'H*1OJ4J ,UI_R1^,@K?\"J+(M8*=^##P2NP6+A\D:?%^XP7X@29QS1
P/+K?N4E$R_H\ GCE7"J3B\T/>2.'6\7G&2LU0,H"#Q^R?[VGH3U6U'+T-WIK,4&/
P^6RM9R\;$5-ME[%)_>6SVIFYEY3Y;VIT050Q]3,E(!I9.4)6 >WY]^KY,(;W9?F 
P96YN42=Q46IL^*7?%G++LR8^.DPK\26%.E0D5K8IK#2VW^;,V2PD4)BNYXXJ^C-\
PC4T0]W'9+]K\T%KJQDEA?)I?B:OEH9@RPG&$1POZ6U8.P0>@K_L<T,YP!3Y-%0B5
P?SW?K OZDR'?PBU'.*[&&G8=ZU.R=X65"T#4M70,CAD4>J8BVKO"S.4]>E>7'[MD
P:$/!Z$A2C-<.SH?>%'R22C?!('\O-:BM[A]R:I=#(EBQK477/P7)P85)WQN@Z![[
PH*YW' $]=5$THGN:'?V4);S>#<5U0@59,NS&&TL$/D@@PP@>NL)J[7H84*,VC6ID
PC"[,J,4X@\$[SG\#;6ZWH'!<]X8GG0"E5031)GN8TY><SICRAIEG#P?&+L>&?=O+
PPT@ 91RF0NJH@,^.,%[<]]*,WXA:]"GK!HU$&O%>I@MLSA=?G_D2IXY35U31L:"A
PY$'->%4T,85_3$NUKLF90$. O"AEC=C##@?-ATQA-D.GQ,(D$S"6'SF?:C_:35#Y
P07Y*$S%N:T^C\FHQ,@YUI/-7V8]IN4-S0Q(3U4 5R)M_;?<@5")0C78LWHY4FGWF
P&1!C$ \@DOZ;-O#0IEY!K1-L6& =.&X#M1^J;MJXB^G89@E@04=T4::58X62:OY"
PN@D!3;)O>IDS,W&O8-*^115$;45@F?-!:]F22(>! ??Y6"TYX??=#5.#LT:!D^]>
P?.\7'@?24/U73X4EB8<\<DND\P'*Q/U)5B9OIXE>NW:')\ZME5 M3UK(B6A 8=O!
P",T#@= 2W"(%ZT7JYR%4OB&1O"1/O8$5)?KJ(#BV6\/?(^E3*/;C)"A]"O!O-_:C
P?&LW#FWD8_;7KR;[GR1LXAC36)4V,7HC=5BT]\%BIZ6DF(BHCK7:0I1AS38'IWBQ
P]HY).WTTPX&8C*,(W"^*]>C0,V18N]8%+B/IVX;<ZR?%,"W=)LQ9OD+J7M(0:P:L
P59?+4R_.")ZU#FX/E(]T(JI!0JW:?4P*3V8*JQRP><"9?=3V 7)-P;&IJ K<0L1K
P!Q&?^_P71^/OIW0-P"80X'O)#+\0EI +%'=L7ZV-G_Y*=OL"W AX5XVSC,DC0,_Y
PXL'8OY[KIIRE+;4EM!4UTSC@,9V6(]->7^U!NNEWFPC[.Y,\BKB631E,.L9[R0?0
PT%V)W[B89$6N,?PQ_5*2(:<+VS+I.I]D#B\GMYUY2-D$>4P1E$:-99V#X\IT%ESM
P^HP#/PP$"BD1BHY&$\6A".OOY8;\[B1)2O+X8<?OCT+!.MLJ"^?GLSLY,*O/ZN[-
P6&:N3? &(*"!LQXO[[&.>8[=5PA/"2W7\*'6/,Y[/!D>DT;:-2,(Y$Y-5.\$NP<'
P2M5BD:EL,X.R2K;QY0OE)1I%)Q5AURK!'BG>2.]R;1UW/7SNRSVR\2IF?XWM7M>_
P2?C&S"@NH6:3K'4A. 4Y_''!0?3*)<^85%/;NWM6MO0RP &.3$T]&2VO<8ZKQMUZ
P%SNSEV"M2O+\HU',A>B<C D(Y(^B='Z'?6;M#36<'E#=_T:'^AY8&60]NQ.F>1UI
P&X<2W@:!C19,0+,'#69M0BQ4)M6#YL;;4C< 0AL?>A., F[=2?@:[K44H*;B%8WD
PNBJ0'@' 0X(E;^H45[I(.XPV4JH_%MTG&0CWN605\SLZ<N$L17PAFSV'051P H&9
P"Z5[W(.D^V!%LN, ?_/N?2BP2^.&% QHHI$]N,;3>P.=3J[Z>Z=?-^ Q<(S[N#@H
P0)%>9.(G,$\NA>4QR$%;?"Q=@40:'\-X&$%7RM,_Q";7_7$=>!P4#+[8)(),U[*W
POX8B0TR/^\_2\XA=AO(H.?CP#W%/;(6#R;3>+7V^UDDT J!FC9N%9;L_/^U-_=>0
PM>F?IT4V%E4SIF.23>^ +%1AN_:2/_-B.!7QB97 EE_W-@4#)C4BY[6A'$J=V6IF
P=ILIEII*/5[;+F6TMBN[.L&6AF($H%$^9E5\WQ3>>M->=HNK8P5R6ZS#MA#\UGR8
PRS?831=,$'YASMU7G$_2G%+?&4_BBMN/NX\BJ)<71\PBKH=,9<LTVM>EW15&@?/_
PV;!/+BO>DDPS'&QF2=WA#:HR81Y '^\PR:$B$E_/\GAE@C])P$$^J3=#A@ :F' 3
P@E491@"Q+GCNKMAH!5,;X-H#L<$-7$YN.++PFO4$D#F;]/I(M*-2KN0(P&Z9"Q1%
PRL53(3SJM@1+) B)JMG(:TA9774E'M(0S!A /C/:5>&9C2WUX?]4Q#$)8!\U^K=E
P-@KW6@7A0]!6P7TOW&W-&2_MY31^^SD?\O,C3<I\$&-U^AY^#.EP?\XE(X>*,HP\
P6,Z467!M?J/":I8,I)]%CNO;I1 ^#$*N@.X&?-27C.QI=E74=8)-<I,,IS/IN030
P!JS*V<UVHH3HVNF= BZZGYXH-2PXB)/DTOQU7G&3RG:E<U+_X9/F.:LK3)V<G%-]
PYIT):3-S^N1ZHM*GN.*%EJ>Z#XF]1N_ZL@?]M!'/D>^[NF,]GTS_W!&N_>N1J*WW
PP84-Y9:)JBZ^Q*8;6;1<.T <A9?.(:-HI,XWW8'*I89MCTD8*-(%NE^)G)[F%%;)
POMDQM(A6WVVJ) TL1AZ5U+0'$.'C1%M:A=;J%BXOQPN"0Z:[<#M#C%BLGIM3S<7 
P4)SSO![*#O&JM\&LM[BZ!TO#HWOS[7&:D<Q6@Y]*/-LW]/.!9IJJM@6SZAK>(ST^
PGK<XY\"E+K<;*:L1RE?S1P#?9X^BZYKYRF);?4OC/VL)CW*86\%Q,5"FH]@ _?=8
P\$BP:18QOJS301B,>Y<MJ08K"ESI-K*U561L5FYS?9<47EPRPU2.( =?,V.PNJ?"
PG+>5Q&M[G9)BL==(31@G'46K4%? R',V@SM=ZJ=B3ZB_AD)-X#6]2-B'Z"9;>+N4
P'. EBJ&^A"N);#(O@?LW<)'ZUVGCTY/CBR*V$)KNI5MK@"B'+^H%#/+ZQ#Q.,O/7
P3]G6<_Z75Y,N4KZ,0DINS ?\CS$^%X>WQR^%\#JY#/" -.VJ03?K*X(R@W?!K05T
PT-LGO?RY;39G+I35#"WQ&O+$(]$1X(9&L82+$B3D4F-XS"@PFVATHY86,.$T9GD(
P5<*/>[*B^L'?/=IE0C(HN03BQ4I?5,;>%E@&)=1?C-*(ODQO4A-YY%3_J1'9#[RV
P\Q5T6J*)T=R-F_H[4/6?@"/##[018VZJY_7B\RB"2^ MB3@-8%<;;RY16>+C6'AM
P?^&9_%M)(A),/3NJ=KG*E^R6GD-48GRSKHK2Z]5-L*6S^K$)!8X8[MPC?I'_3.]B
P-];/?(JJ!]A&&<FY,?@_9GI9AQ<F2@#].?@J1_I!0VFH\%['*&$O:J-L>:DZ^7,(
PC^K]2<-KER?E[YG%1OB)-@D6I756D)/CRX>-UYJ+-AZ%#@ N?6I"+892_TUZ;9[J
P?ZK4P+X>-N&,>_?*LRL<*7>+M/8[8>IB6W,>Z(=Q.YE<"45V?\AV1CH:R4=QZD(L
PD32$LS99OW[5Z[J5HEC$+G/8NED"CA,&-JWH<$CXJ " I*[@5]!KDO'S<> V;D@U
P@N;%.K%<Q?#L! ,"PAI.BMZ#A7C\QE7^7>7/Z0($TZM3$>YLBZE@":3PX20VTH+M
PPAY[K*_)B!0^-LX(O7%"R#\N(<!0&@""HKW;HI_\UO\+D:VQA M<.I(RTD/L2S$@
`endprotected128

