// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Guard to prevent multiple inclusions
`protected128
PA-_/Q@:&[',;ICJ[?.MZSX,/$DE?VGS(&S14^N6OP%NS67Y+OTN2PJ3BC7N[0U#J
PO,YH".^I'M:[QN_[M))9FFXK8(O<>3&QOJO-&L+]R9XI[4XXTB[S_[+K %F,5\KL
P<MSLC)#'>5R.:#NGNLE6V?4K@92 ^Y>U +;)P':[0.53*)2S>V $R9'LH?SP*)R0
PNS2##ZHGF ^<M@@%3).MD-5^JF0$A/$[N5A"-E8%EC&/_X5DEG9'RN:F[QAU;W4T
PF!ZS61P0NFUK=1 UQDA*LQH0"&]7/8OTA+7\4HURB9?'Q>@)=$E?L%UO#EDHW!OE
PCOW*N_842%!C/8EGEBF8<XPDA[(U+V#K1,BT/*+0=[HHT1%]* IB:\F06.P6^'.<
P#G16:+<J1-=FO8IL4Q(QA$8&?-4@,=PR:+;F1Z?92R\@"D@Z'H]]%< <G423,N-&
PQ]ZFO3_B $Z7K0YM:]G+?0W^E"OH4Q5K9)J%BS?9$4D!/7">O!S1K1NCT\+:Z<*(
PTG9O\^Y-6EL,0"**6>^X+M9-WPAGC[%)]Q["4@J4OGU"3.';^?<Z,D_$JX7 Q#U0
PPF3*#H'<)7NU6#>/T?T)_9R$R@ZC-D_QS2BGH'@L,NV-(!&<SV,WC(K5 HZ8UQAH
P1_^DUI(6AQZ@'&WF'Z($7II3OV1L0IL!1EL,,IPV#>G 3F_ZP9&:?'U4C%];53?A
P$7FG>#7H^W78N0MK%M0D%J*"BSIPGMN;DT"C0P/XZX3 :_;[TTR=X=T@F14@Q:&'
P;%O'0"_0IVQE#SQ_@,I4^>'8:T(^\PL6 6V784T=2I++)E<Q"HH^QDT9L'E29[&\
PG2[7YV?-"0%],-$'Q7\VU6R]?@4&>)?/$"KNYC@Y5.O5Z/1!BP%@&KWUZ"R'+!&V
P05181^+.1:-I?HVD1I!*-L]#YG0 )A%F7AH-@IP<-<>ZCPF8,#P4$3S[[ =*A0['
PVG! 1W8V]RHEL4&A9RUIHMZ;"YEUI[H;8V62-$ZB=><;JMQ(WLQ3WS>FJ$1ZLN(-
PAT#F$P&%0UF,TV#3'=P>WWLKLB.[[TQM"P%G87+\&)@M,<Q#PN@X=+^FP1$RRJK"
P8*H!EOW/8CH344*<6T>9A-B2QX@[>7I66E0MLE=VN]E<U5$C+?_8OU._L>J@N2QZ
P0TT()V 162CZEWTUK1N]WQA#;P5R%XAQ%[^M41N*M+;!JT#;8-LT.]7[,."M@P C
PSI(+ @\KW9289XQ>L_-MIIF6,3WYA$3#/\]]S9%>,\2]6K0@[X*.S;,3<2OYWNN:
P-W3;_K@-L*OS1AOC_=I03TX*B"0TAQR6IJDZ(!J1[(.0>NG6F<^ DRR8/?SRT^<4
P_/VB?4W!_DV/AQ2V#D #'I>G4GM6)H8W4((35+PU'LV*QP+A<_USJC#C^):$CT2K
PR"+A?HQDM2KJB8HT<)*U@-+ZM:N?DV:A(]$-!P@VQ=MY>NR;)>JC<5.O[IUL\=5@
P&TK9[@&.S)!K.9R67,Z9T3#=XE'.L5W"LSHG6W+&R_N;7,1\>_I.>,IS:_,H!'+F
P'&F1Q,Z#&Q'YFA%JTD>J^D2:?4318D MKA.U>[U@,#4,!IHZ+?@7QXV+4#1A?$8%
PK&4C-Y575R+D5J>&^'!;TRY?W&+U3YRO2E4&,^];9G"QE\?S)U^O)/KS@+KWL:1F
PQVG<(FBQ^#DL"\28)\X"D\NI?1!5"B>?PO.HH8=;%>OB;%*#5G5:0?Y(YIHG'2I'
P8 ,O?.FE+#CR+G:K29%^64>*.TU.1)L6=#SI'ZIGN]EFI])\7=5+);I84/OGCUPX
P>:HJBD6%<NE0T%KL$8K^%NH&1)%; 5Y9=^;XT=. @T.Q(>"@2E7,+\</8^NL6D>4
P)7[0T^"69BHH!.[H2\6AN4E6(M050TYT=7 S=_J34*HI$G-FXA"+ABV0[,6-,-M#
PJ06,GD_B^]A\CF"<D;Z'%!2LBX@+4.K >K045WKA7B#FD9R<M1^1%C\B7:OYG9QG
P8BYF/VA%\N%;V*^XP5-#?;ZGX8 %&'&.QP##K1(=0(_,AEO#-P1^=.;.C93UT5JJ
P+TF<,#I= 3-=UHWP@&%AFURD!NMN=18B/2? YH26;&3$4B#'G3<QN("Q6I2+RT@>
P=2J'J>T?:0)RR"S5KD0I(^"_61.9NZZ?LQAZ 0^V$GS)&Z$:7W]48MZYN;6PUM?*
P*\&3UYI4)XT@LDWMS*D?<G]Y9?#1651;K_Y"XLN0W^C,6>B78FC)T\?P!\D:> #M
P[J/N*S[U@-Y[$7MC;K_M\W[# YQ2:;MN/OHDSH^V,=CJ+>(4MY8<"W#9X$$31R27
P-1E\@AKBS,L3YE$UY[OP5ICP%D13GL(;^"<9!NS,'XLJ)NRW7;W@I4K8/!F]7XMG
PGH1T98:0WB[T7#_]&,RA5N&23"'B##'LABBK51<5?_[D%@FIZSJ;3-M'2(5 Z.&9
PR&GSS2B^PIU7YT$\8Q@<]HR\H5>(+<1999G+3R<@G_AU<_K>[6\/QZ;#S8O(BS"U
PJM@G9(86Z8N+!/^05$QF:\?MHX#P&Q=/J"-;Q4W>=\KM_8KQX8W5$W;?)CK7D"/#
PTV V+)\UVKXO2B^AT"&Q0TRP][&T7]0\X(K+T_IRBUUFW"1X@-S[8?<1.IM&\'8_
P-CADX1"$\=@,^I:G9%0X.!-MM^6HXJ/I+=G ?_2Y5-E 1'N_$'L,P!X?0C(015[2
P@7!4"*:A'ZW_ %6$H#H3/D]""\1ZP[[^@3Z,#C<*>2:M[3[D(AH5U-P0V@8$6>^$
PBTZ<=O)MVWMV.2NK@)^LZF'#KZE%+BD?_&[DG:T%M3]324N,'Q81?,I3K_7.NI$4
P77FS^FV%LM&\@H&9?SGQ> 5!(W/^1K\Y,--NZ%4AEKJ6\=B_YMUEW+S^Q7_#1["-
PE$C31O,55O_7>P\Q,7)KK-MN;H?_/^I3^3((U"Q(+4!T,W'CB=ASOT?LRUB6D6U&
P';D,T3K\*/PP\X3&!&GIQ-:WWT^84*M1/M8R))/XW,G6JNM@$8__^*/JYZ=CRU&!
PC(+CZ(FJX;C]FUO<E:9T0%7!N:-4Q>S^3$$BNAN/M]M\7[,'ZR_"I7C/B1Y-E\Q4
P=G<#9<_/>&%+VZ9(K1;$\0.2E,61MK1C<0P7X@1,,W9^..)W'9E&;&-H*X1"'^K6
PK!I"OP:\")71+B'XG,JW,34VZ9!W,7<KOS#!8>G<)WH(7@CU]6U[<05J=[(FB:U/
P,][X%/*21*MA+%QQ$DCAR*&M!%%71;+M>O5 6:R2C!=ZOF)$U:@*/,56R@>G,W$H
P8#?0"/0T9I^1;</M5 \N H^JYNZC]1C$I8+OHKH'++0@;*"/H2O-)!D](=,9(^+2
PV7 08]WS8C"Q\^%)=Z:*(M?SNDM552&P7!+Q4&8D [[1:K9V&9<Q]X,I)6]$@LV0
P)ZI<6?Q9=7[1FQ52]V8),Z^+Z\1;BE(Q#4C2/OA,B"UEPOFHJ1<,"'_[8Z @7@#6
PM4NTJ@F?7V^"")/9JDM1=T<!7COS3%9IAM11]:#G#T"Z?CNZU_]WSN8!X0O7_L!.
PLMKD70SR/\0BGPS&-$R5&>C$[S"5B XOL.=!2A_M*\W70OT@Z=[I7<5W.#F:2.4=
P(*E.5] 2&+!,6YIUFVQEAFIE4IJK<C(#$O\G7J:$O$C+/>802C;1(\4C#$((S61;
P&:/F7ZMJ @5NIJAH 9BVII!^ 1';P%50'*X,  _C'&F(% =%6^MBTT2PU0"1$$@&
PWERW]8/J=8S\DS9DMPQ9_2SQ=ZPJ$I6_ED%X6$6Z%ALO[JH/@J#JJ/T@FCZ\ *M-
PYY_!$[0@[+N;\0Y?G"455\KHJXS(C:RZW6^F=,"J<;^XJ:G?I!#GS1F"&T,'VZ7]
PC&CGOIK6/$VB1[U'67T9;*#V#GS.NRBZ>'."F'16!B>#TVC.!+WKTQ,164'$DXBR
P ?L,]9FA8T ]C:H)&-''L%L/5:"1/>R?3PTSMR[I\(_"6*CWT>OIU@H"Q: M0/K+
P.GWPZBT,\LYN3UR5XQV@4?*1$E"7#7!8HVE!(PGTJPF@"PRK<%U8"4EK-3ZD /D=
P4-5>W>5C=8M( GO*SQ.PE:!?2IZ$X@N4E<99\JU]WX'N^AW5+&?AJ&!Q,O^1R=<U
PD34QWEEMJ8NC:4#Z=M1ZTS!4GWAS@PY_V*:FEF8 _$VSM'72#@\I%RT,X^\,F0GH
P>*?,*K/W>\\S43W X:O*%2FZM7!WT*"XP7WPR?&O97/%OBP$1O;8_^BS9-%^*<[M
PK7^5\/1\%BP^Y91N;S^\OSB>*SKKB D57Y899D!,*RK@9[4$]L;V4.$8X5>,21GY
P:)H3XZ'1KP.) O\S'0F&%TOV.('>$^>]AK]9Q%I.C;?%_RYR-LE_>76V0;($*U1(
P/1>U:V'K5&D-=FDI5VP(4O+GH37O51'!.!3NA2A?;<%V!\FO?3RQ]QS?@5:8AB=3
P3F5?]988A#VF33YW+)%[+JEILO2G34%$A7Q((QKXS\OUTZWU2J*A8\Z=VN&'K*^_
PC4!W^J9LL3PP'^!EMV5&B*X\XNDCG<20XN$#0G#Z5AP&KF_,8T/=^>@LO]#:X^=X
PLX/R1W0/L'2JW%GTQ(PGBL=RCA@NQ1*RP+D1[>[%4<6KZE[IN%(]FC'K$!T*)&PQ
P+Y;'>WX6:LURP#O5%\\)"K%*C\"$Z5"5.JWU5(6@#-D%2W\W^KOK/9FRM7MIN0D*
P48L!"<C L'29S.'K ^JEG-;KH^7%.5L8RGDS!UFAZ#!4O*%@!NS5T<2*$_Q[U$ E
PZ4W^ >Q7<U*LE+]JS'E@^;ARB-FN+)1",2<*V86Z%.D%GQ6@C]"@:DR$*[7&5HS"
P1\ 4-"[0+8& \S_=@-$N1F[43)(OM_1<&Z;?SH)2IMN3,"-@62W&GWI>).9E#! ?
P._FMJ/M1+1I-9.H6=)? J*0 :"C!-M"-SK+8"8?ZAOME5U,;$Z;L]L<'<26-$VTZ
PS)S.PEZ+)EURG&]3R0_7G&4")&2(YNLHW"-CU,(0/$GJD'2+G?4C&C%LL\FNS+C%
PE5(&1!4)W89P7TEX[F-I"\4K:2IBW$L]FKY#0A:YHI%/;2,49O]W+]S/2WU*G_D^
P9QL^9JZ))&[]^8#O.^EF,O 'P<Q_K@Z79 P8T3AJ)#?(M"AN.*;7E*\[3_02?$C1
PLHZ/*_/)=76 M0D#R[](.-,CI5&]MDR2=+L?B"K*?$4*5?AG9[T)PC!PYL]"J">*
P_+\Q68902TRZ1#XOU?QY];]$U_8)'G6ZVMAV[A)'&A)M["$H60G,RRIO?1!R^ ;$
PP,4_Q:\X.&&'9R+OQ8Q-FW@$PKSVXK%I=\P5Y>F'0"3KB]W**)0;D.T[F?&H^CBO
P"JL=$SZN*,'48\&ONJ5SFM5LN *IGR&2"(^6QQ9D;Z,<D/KHT)8ZDQIJ:>FQ15V&
P+W1%V(@2*IXRIM.F#EA1/A)*\7JS)DX>$?PW*%%,) #-"H=U1S"Z#(R+N'VJT42G
PZ< :!S:/YF _,Q>D0D?@=XMW;!03 LAPP95 %%XI-QBBQ.K1#$X4?NN>LO4AL*Y0
PM_PGD]>/_J_TNH,'S,]T(HS\&I<+ZBOYV[$=\_=)9!UGU$D="'">3F-N9,G>P''8
P($;ZX$/P< #1B9TLWGM<)'=UY\X;...":(R$'M>H_"&>.FU@LAQTDW+5Z)%K2K:&
PL7"I_Y<&^&WY45/>#?Y,P._V02E.$(H(6+248")@FWB61$JU=>T5.@["(\.,C, I
P7KD?BYCIBG77OHOFN09\Z X^U))@A+0&]1/A!):!,#^PBJ6QE;)"O])GTQ7#D]Y8
P^C(,B>)3".U6\*.0]4K(#G=JZF>$;LHU]" N6"-85H720J^3.GWS84*EGI-'? '"
PRUJA9( $#0Q#6&K]VGSL3<Z$,-\>8O#70#_=_77&(HCZH5N,YE5.J]1KI)215911
P*5(T'$*P$#$D $P&K>!OU'>> G(AVH>J3 V#H26/?YQK]-(RO:B5W&#-E> @R;R&
P;SHO"A7MGO1FO@>/Q%I9W#_.%U8P [E$-NK/U)BXQ6QU?X,T I>[IL2 ;&>8)C61
P4\OU670@;&WPZL0NS#$IHW?H%K)DG,KLKUM( /X@\QB.Y'!LX2F_M4:O/5/NZ39_
P40-?YO$5AS IHIHW"J#V!Q!NM_WI7W8DSI\-?=_KQN='M$GS.O^!2A60O4@H3V2.
P$VTMKIWH6XCKX58H *$:N]MTOHF1-EY]-4!6=&_-&NI@'=&1R6(($;JL5/O>1RO)
P\K7+%Z( L/9&FUVYVW(*,$:_C$, "Y=OB8\;J[;8U-TR]JLFI-WY??[:+BR-.U7,
P2;LA)S56B(1!?_=35BZK!&,R;W6C 3P+JN( OK@@_E3%> HHKNHU &_!8U)45ZZ,
P9</<0YV"*:D:S;/\JGDHWS*.[OKL(>W&;!$,%<1BR$;YJ-R1>0+1T77VNZ6O.D"7
P_IM*AQ=U<>2]+&KE&->B34KQ];%T_65+1K[73@JD$*9PZ-LGY3[O/M.8\5GRTW%%
PF4ZE<9UK-%Y;C!?"=+6S$VHS-['K?>!HK3"BY3AN,/=U3"Z]T2:X?JS,;"Y&A:C_
P. OQKBSG%-/&*X])(K*8TXJS1$#V<.8 SI6'P:$HFW9_2@5@W [KBBS7@ :L@P#4
PKD>RO.+R&F*P'QI]+6<YR_3A/>; TM7S,HJ 4BW1SOF)0E,KC:W-:>CF)K!-9%DA
PQE//SD$)9)-NPM\'"9:V_Z=WO27"Q N8/:P)4W<)9!.Q=$*9^83;G_PN=SVJ_\$#
P>%^WPH/8S'(J_8TJYDKG?P!F1CSS;\&BV%H_E/M<?'G!N#/VP.UZJ)!P;SR-^T;H
P2O;50?8<S?82Y]. HTC3:DS:Z4XE.$-+1,_/!@N<J_KT4\+DAF\JF24/O!'VFE=]
PMY@X1,G=53N2HW+.^* 96SDGW$TM)$@)]Z']1HJ_T(E\2P^80X(GA[5E_#<GN0QO
PQD,%5G,26*8+ ;\-8H<EZML1@ZPCAP?63C\<2^1N]DG P;[0<DBE_WR:W8>C =/8
PK4:V5S7S64/>\)3Y%H@>'C-&.WY8[$5>!.@<(0IDC[KQX&+DHFRZ:3X.2-;Q49F"
P<(-];D6)I$SH;K*Q=AGRY,$ &$?".V6_U#VE3YT!!JVH"]@QW$ 6^9?$Q0@&&>0"
PKL(S_J=&4[A"-YW:6G&Q8>L8"XTRDY]7DM<&]&[CV9 S[2T>;T7 <G92-"WIWZ")
P5-MNVE78\#Q$5)50A3A/J>T)E_C!X7SH!8XYRG\#3ULADVL8QY;QLB43#4<-<B:Z
PC-P)#T#F. [,]4J@L'[7L9IJW5U_8!$C\<O.V2$Y[TM^2!CREP7XE^X?$6":SJ4<
P/FM8.H_?LEG2$JI0OPWD#,]'=M3AL+6-XP<MP;(W($8[)^.5G(:2;6XD.PSFO=XN
P[BX"'W8RSU6&#1MF?A*2GRG)?;%C5Q0P-+X^_FMN!1<!@3OK[[@<&.GD@<&[PNQF
PV?1!PNP5\$]7"@04H=A@%69P-([F9C1+N#F[_<T+  I3:)VV@FIC4OH*.7/%T"*,
PBH4YGUM6IYFZSC+<U^TCUG9.620;YC/RH!*V-;]%6Q^#R$(0^RV_0M5U1C'A+"@"
PIL!R;7Z8N:8"2>.PVW;&AQXN*$@ET<@.*=[*7GJ@98FE,+[>=9V PX;.-G@>LH4=
PV)D4-&V/BOE[<2$(ZL[< PNP*"VXJ]_R)5/_EA$4AIH/N2F@OOSS]1? DM^ZW^&7
PGSWP1U_P$ 9 P_I6\A@IS>IZ^%-9G^\^61N?(Q^8/KE?5_>P'G5X$D:E&+U/16Z9
P'?UD)$&'BCIO9M%A@(Q4/:>2A"N_?61-)V9/W+KJ^M*YOS(AG/VF[9*G)EF8XG!2
PBTQ1OZ\ )*#)^J6;$G['E76L?\X#*@FMNY'H]XA$Z4)7U=\[Z+X.%)I"V+-3O!\2
PH+.!7[O#F$5A.PI=JDAEGDVM[4*/>I:17L!JC3S,,33HI\\>CG2!47(0S?T R\PR
P/M@[O"V-B+DEC>5;(G7PM,@O]E&R?>CDB!IL>?R^<#FMR]!(&MVF'\ZR;!@0L"WQ
PL"'K!^OGM;&\'(.XNCX1NM:;KM(36UROD'1RS[^*RN9QJ@R'XNT^@@Z5H/$8HFSQ
PXQ7IM]B ,19Y5$W9*2L#Y?&'+-3?DRWWA&IH0%(E-*6UA:% )I]DX3UUC,W4F3B:
P*6=Y?K>>X\>S'-5-"?UAF\K"Z0@S+_82)GCD"9D],T?N JO[I$=HYCF#VX5/HBY0
PI6C-HM.[(SL8S54%'&4"4J.#Q<105$1XG%=I#685Q,F !\YDAV^4\FP.]#G.6<4S
PW9I\#$]OGF7FE>]"=X2>_0-SAM".$T5.G7\MJ>W!@6MK2H$"++\T-[%WH4.]I]H\
P966%<I5>33+_A#3G5+UF"Q2R7>)_LSF"6IMV_&XPG>/1HMQGOE0B,TG9=_&I)2$C
P!/GM'KP.L,]3[2X 8,PD=+]8?"RXZNAI*@RL*YFQ:#X]7/"L0^+/6K]G-"[5G,ZM
PY6<AU4OB1ELS_^SP5)5@YGJVN;$@PF5\V+3J@4#PA"X8'7EQK@Q]@G?ZKL!">^1$
P@/CB64=@XN^=X&!U15BL$+N%_NQFBM>79-<I3ZV,A<+EWJZ8A,G*#SFP3)Q?(753
PR^0*:C7*+G,;JL; 7[B)>!/N;.RHNJ7LYU S253Q7^62:":062[8D8G(%]%G/;.K
PR(%=DDC]43AV-XR,!#@)H,+QJ[S98FZ:>T,/\'&/,AJJS-FZJD++(E ?:^5.!,@%
P<."]=\WUHTN7/--LA!1-?=5TW,]17)F.E[\P-HY5AM;^/]\OZ*$"DA7=(^.?V2>;
PUQRH5VK_ ,7\0XJ8*Q?[UW/2D>:%S8,NA.R9 4#@PS-JF?^;!U:!I/()'& @.OB&
PRHOM7U&!VT53HIN.B+<H?&&^L;+3'U,:.)N7D:7<UPN@P&IB!QPV0U2QPP&BW-+L
PZ@Y_C<KKPI[]&%)?2X$B"%/O-6P/<_T^<S3$)6:)]'/*"2JT9[M."\8-.LG/-M14
PG1;)!,IHWFIXP:3EYRO^S.<#WUH5>.N)9_MY+8KDTVA /)T_E"*XQ2A[U*^0A#*5
P$RP^NC1?9$F%KJ_U;ZALZT3MGC$I4_X>7F-5-L(Z(G-:V27M[V$!D[C%A/Z/JAGX
PE&TA\D&'*.MZC133,' $:2910>0+EI7P[W$3U)]="7$IV;<&?C2'9LW2I>CZ>B',
PU88QX[YH364'W$5C9P)&*-MEQ&S6GNO:Y321CXK[6;$S$'?(#T?AP1&&+%2 &]YO
P83N\'U?PUV"='4_XG41BIQ5[]]NV1'F-#37JG.B/ESFEI_LY.'XT_#-;+(3=:\SV
P[#XS(;4^65#%V[9KN4I8;?(L*_<D*K"J6R5PCDUB'_ETS==SJEL%L+8]6]4[.V/F
P^L,Z(S_$<?-2-;_*3"#CA33S.^8-B*NFB%X>8Z!PUP3 J,A5%X7W-URLDQ8. @H/
P'%Z4D%D#Z?5G8YB ]ME0!!9D \9E::*MM:Y9&3.@J""YC5;6S8 3@0TS0K8+CZ^D
P>@+??N!L@XX-8.<YPK$N.K,()]B=%E]G NRV[.?MJ'@)\\'P_==LL9-VJ+Z/U-PO
PZDRI+DX]>-:OC,88_E:42D?I%@+D&WN<,7##)B5HRPBULH#&:5314.F4$'8MI;U6
PBD1OWPY@39XT>5.RSA:]3.<M$)8#&;FV4Z.S".-@XD6J8L!!N6Y9UX^!$,?):G;$
P7R?E%PU9LJD[?A'*4ML7>#4S'Y>\N0*'(/Z,DWZ- ONZ"J4!FLZH>LYL42@)QIWN
P#*6 G=ZK/4YG8D6D?%T5?@BERT;VB9X;EB'W9'Z<NB7K..G>4WC05N,C4\*[/AS]
PG#SS(K@+2R9$\B)K@14]^G3GD1H<&PDMN>3.DD? UG'L:?@^'Q)53RE.#$0D.'!V
P-JDID3^#]5[(QV)0 A+$AU8I;A,A*&I>GS;D*RJXV%3%O!.FB6&F)3"QSNL$MB62
PD6'FDNG;GC$,M^RIKWR_Y@DL+F?MKWT:7FFJFGY_Q10J^TJF2E, PFM\8?K&>0*V
P/-X';&&,X0WPHE7!V!IKL;2>&A<4 _$HG\WKFTZ79?PMR^6!1Z8Y/1&HJ4-_2D):
P<-@?VRV5#8R8]90:]U.3$3^WH;5&1+SF)>_$-!)39/S:LR/I,,J5RF34(3CFFI;:
PNB- HVT03Q!$[\(HP9"\B5A6O4VK TO8G<BP!I$T \#BC/R=<$"MD9D=0Q0N...@
PY@4:PU+$[R0KM(?#Q*LE>1]<=ZQ40S)_'Y@"C&;V']0T<L2ZS%NM\4)0;]RKH#.T
PA^1D&=R972[3-G_Q2()<-D4>DJ$OY+Q>AMZA_O4J%> ([Q42')K4TSB00Y?OE?:+
P-!/E 34,UDM-T76\GO?8EAE%9.[5D$$7$R*T6V7GML<P!M2@(*H7V<P*6W# S\[M
P5*Y"VH P:TA(S:Q],J(I[8"8,J0Z^67$J[B+%]7!!98]_8$H55@1,_O\79)1[P]L
P\9)VG=C?Y6:W0!P;+LJE GP]"OV*E^ O9JVBE]K/1S:B]2PAZV-^TW$)[#M#O()0
PBU@UNNI;([Z0C90\WV:5XXPZHWUJA@V "#1K@RCV*$NE?<[2L^NF),R+9*%YB _"
PH\8,6-@ZQX$?>E$VMVA8A@#\B1V^UU>V NL]J]='EL+HR;04\N\/S JL\8\AS='E
PUUQ):6V;V;\RUF<N!8,^LU42VC.JZP#>(SD6*F/QVIB^^5K>=\UXY>OM+W4&B^Y0
P%?0%219BG-=KCN=H=J=#T\(URZ\I:O1$$/3L=-EZYXQAM,V_2#FU'J^V^;6 >*-7
P>+S;3;QDVZ*_8S0WRRGR!(8L3ULU&5@'QUOL;E-!A-MF"B^ '_)N(M5\KI.8CI"R
P<8N3+WOFS%8<Y>H:H6/U-AY4%#G$\*H'Y])&S5I%.7\>[7I/3[.=+C0A15'[0<9U
PV(D[-3>\L.?0-(L"<SN4<>[H2J?$JB[&XFBK&<=4=J-@$-&B'>[;&C:^8A 5 A'^
PH< CW:;'$"!IM75"LW\M*W*L90+2YD)]5URLN$+6#NJ>19I2[^!B99A\O!TK_9<%
P;(G4*;\L(DD&<XDEYEX7;Y[\CP';H('J]^_BG<!R;R4#WID%E:"E -$=CIVPF+0\
P-T23LZ98B;;&:M#W;]U<@(6#K77N H;BT<ORTKJ'\6C+'D*^=O>E+YKEEJ-\1S$ 
P/F08WRV!8O;U1^Z54VU*Y#^F8X&RXWBETF$P*%Z7L/A],L->HQ[]\U*C5?QD2=Z7
P(<IG:_&N<<,1=4%Y%UU\!.7B@6PR7=?MFL=:0'I+0>"(AR?;@"G:?G(#&R.!#FX9
P$15,_U21ZM=:E N%9S].FG,0YSK(,9V+^7RHF(=@@L7RBV V&&9^72F!D45VYZ_M
P B7"F\I@!+QZB;[?RJA6(/1#6>/DQ @#UY_&XD7^J3Z)TI#P^^YGLF)#^>W>B_/'
PB9EF2C7#7?^)IL$[@<'DK&"E_+?G#X]0OV7LP'G>#5&7?^B;[ZOQU%'! $)?;M99
P).D3GHAU@K?)ZS-C?>P819M3B+2P.E$G(;.9)&>FJ,6,]#%K7XP^;7:D46(U7X/.
PSJ-(= D4BA(TQSWO_@3VC!B'AX;":)&T.++]EH4J683-_L."1-):$KDCMV+49P21
P>?]F978&*L'4V;OK65[/Y)[!X]=6++L\B!0J)4N4.;9IT8UN/P_!2XEV&2O5O15U
PO?H>0:%^PFVGE;K547_PU7Z#L-_\)Z?3/YM6<80F4*3U*X\0I#<8^6=2GE3*N^JT
PDV-3:PH9+L8LGFM_2V@CL26\+Q_8^DM-L0,-^)7)<U&'?\*V*QE4DLTF-T.B%"TW
P5[%OCP1F^2WK1Z<L$9QZA(<P[4S^TD5D##/<V+Y!FY&_&(D:L -=B29T3PO;O7H;
P>#3H5BV CT8P!4JV' Y*\F%"B:R_QB%GG(BPP4BI59X:7Y3&IZIV6-F-O2@%#\7%
PZ4X5ND3Y.-Q!<PN<:^M&M+C\U$QS^\T(,VI;P!LCE!J_3U4-;&_21^%=OAX%XDL0
P?3N:/Y^"2X0B*0S<184U:'WY;J4 'J(S!M-%BU@CX:KR-3\Y?6Q58=FG#!4-X.>K
P]D _F",\%D$^[#?_L5% #R#YS4-_#A5;+8-@1LPENXZ*&+W<"KKAIEQ3V>F1!&#"
P0H$M3@_]T^1F H:SH"U"O'GZ'FMKZ^!+TS:RI$F]Y=GDP:8$7TOW=8&EK2E*-OP$
PSP]/X5MWA3Q.*48Y,T]B$,MEOO%RHX6)0=6.,MSBA.OBJCGB<D^\E?3C1 /%>1;8
P0N$$K36N&$SR>S:ZNQ9:5Y6N+/8)3"!V[&PT''-6H6,<KH;[E:6"K+SOIQ%?K!48
P>1.I+0PEL$EB'O%D)N6#@LPI&I)3/59&Z:OV;XUFUD/F198 &Q/':>Y(V-FI283<
P,K4K4C_TQ],#.#/WPVU,O_*>#R% ]XI-+5E0S;#SW'N'"J*DK7_,7X?C X<-R^G_
P?V60/PN( T4\+,4A$U0,5KJ+B9"(<7B]//0VM2QT[$_0WAG4'1:YA#4X#@P^"B#A
P++G8\,)FUS4I$ZKI] [P,?2PI>X,>DN >@,TW H+0FA,!1;K/K9%- .=-9:AAV#?
P."'5I3Z=YUFT(?D :OC!>DD\?GC.,N)X&PI@^QQUB*._.887[ER:&"<AP!S90"/4
PBBV)LV)4?R(_R;*UUF93IF*;G_#UL$40XR,L##$&F#OZT(?5_H^D_<#GS19O$A J
PUU6*OT-@[LXI#7R4_.6BW%&$2>K(4YMJK(3)]#$V<:FZ./-E>RJ".Y5.L80=2W==
P2FTRIJ'D04F@R6?.RY1IF03P  >ARJUKZ4F5L3^*XCIEBCW&QSQU;1%.L[LUVR6,
P(5\/I*"N1VPDA]/6$0ISZ$X3Y*<VVFJ4Z87GUS>LY5169O</RN*?AN!(H)%:_P$:
PWR5G#6O'2AZ<N35\CZE :5YOZ,9=.<I,N#,]&+BX8W*L*2I=7G+I79:+4<QOZ3JK
P8.PJ5(0*X$:$I2HXVB"B$FYP*]4 &4%Y6R[7 :>53((JJ-^%2<ORWF9&GK@C3,;L
PV[-JT@\$73E5-!$3V9 .:L>VSI"+=GE=>OOK](F@403CC4,;'U@O;YRZL.^HRZLG
P89VS1$3>.S8]UGJ.PO/$-[+4K*V=6CRCMU&9Q[W#,>K!46YVG&LP=GGB+T=O+B7F
PQ WH31D"U]%>N4%.+1WU)V*\4Y>E[X<=[D\[C:3H?)3'6N F?XCV?=M=O+.:'<6R
PAW;XIP>YES>JE+93DF?^9L8SN2;SNQ'7_Q=LEOX_%A+V%T""Y)7[55#T\L(F//[J
PA6P0 <2=T'$W 7F-[__<DZ\N/.5>C*Z*[822E8A-MMW\&0S:@]$/VY(F,[^)=(*Y
P\ ;QWN0FDE8!4#A_6-=\ $L+EIG5LLPT.V&7Q*?XSD%!D-9[(\A*DSW!SC.0H-G3
PET"%>@7R40 &%.:M?9I/[ E$.8.":+K^R5JAW-NFJ96] QK-Y2RT%6:<OEZO$(:#
PF*9,TUR%KEG=A"+8F.(V:PP_?>7YF/E.N*IL "W<,D/?6C ST^5YSZ'0'O]6C6/H
P C8"EM8F^*SHRM)R!4=MW8OL+T-%Y,[P[C#EZY5 >>[&H\1799#=IS],@]L,;4./
P:V<F+<8L*7@$IN=ZRGV_B+>:#4![GS3EK,?5=2FC".P!ROLP$Z)'>A#]Y%+$EX^*
PJEF$-USK4.'NW+[5TP67&>OH67;[BW$R[06G>=R\YH;\=@M<):E[@EQ\4&_?]HOQ
P#LS$KBK1G1YQ*-3H#&FU."*D4S0YK+ @%8"BDI* .6;?N5Q@7_I3*?YZ&7FF:,_+
PA(OV>I4[JDO!OZPL7^\$/%\I 8.&,8-BR!O;W=>*0[<B.7EPO3[.[2)E*I:]L;*F
P\MIVR\IV4-/UQE[-(>NP/:-.4W#B6A4B7?J=!3@Z^W%SN2&<[?]/I0^S.7;&F=E=
PG$Z*CD8 5XV5SL*Z:16B%#R!U8S8:-)2/B7_8[?X6DQ+K>>0W+F<5D;0I6R-603V
PGC\B;:Y8A71\/4%/8CI(2YY*!%=67ZP")*WNGIE\/#Y(I>N2<-!D$)'>+M+C'00/
P/>9-F"Z6[8SOB2_[?J0^>\Z>MO'K:/^]75D$0S.;QZGU4!^VF'73M:$ W)DEFTL7
P*SC+@\MC1W@.78A<K-'W(RRU45#2.O'FWF>N'UHQ9,G<G-:\$#.P_-G65@'O^:=4
P;#;6**V*ZW9D#]8'!H03[N!F!!^$) ]X&@,7Q[";_IWX2J@JAJ!JK_B&U@GG'FEC
P=*O&@^QU:P\46Q.,O1@!<43@'>,D0O?>\LS\2B<C;II1=SML@EASP<Y7(S]($@J 
PVTIC &I:^3L\STVD*6:(NDK[N&:%_3B#08V:%-(]O2L6TRN-:W*!!NA# <84& LS
P&P3G=RQ/;#9P]25:;; LO21SO@U,Y<T).C&10F9\20JL*&TGCBBFN_]O<;_[L 3H
PA ]#3 [^=/O.>8V\SS=^Y=A(-56\$.C3(OU!T<_OA$@.GL<Z3N@^O>&WP#@,EBUR
P.78\G[F+S#\^6))ROAF;Q3FOJ3Y0L=_J]P*G/VRJO9W[R;/D=:>[@0=J9Z+6NI)4
P/NTK0HJEF2('Z*A*KG4/S<Q[&FF4;_'F7& :%<*Q9P3:IL4?N59&Z<JD.A?P<WRI
P CW_J4M,*[^^@[6H9S+Q(LS!>]R<;IS^ RV5N""%ZI$.2S'H-*P,58<]%X1WH[OT
P':FSS[&,#-+LF)DD<05S8P9$Y\)Q3;OW?S6RBQE\R_8V:4D:L?[>7Q\V.K3+ZPL_
P?BP!HK%A^ZZ)G"%$):8LI9XJJT_/?_B1)3\7>T\2#B%HV'-\?X2__$(9BFL\^$JF
PF?;>1)2?P(8T32J/:3D@$/6%4X@3+M6X8R];6O(F.(?T5 ]X%\?L348YZ*Y)C(21
P0X9DX,RUVSA!37 ZUJ1UEP+70A1WS,77AM"&8:EN<MD=PD/*;X&Q4-[%D;&>"$3[
PI?%X3TGTJD/V:X0I/?RH7?ZA@AHJ+35$JF#)#!,/X_X5^T%1_0J8L\7:G+#.O?]W
P%XB?0Y*Y;>(';GG\3]U$/7JK<>8:@9Z/6.8Q) H \LN^;6+;,'^];A[ MZBQE+==
PFZS"<T9N;#"CV?U'D'ETOKMWXH(RN6(;!-S9,%J#7J501SOZ8SNPC41S!8TMM(,;
P),DF^1794CYT]>WAHZKBVQ-"")Q^S>MP CU\9))J(4\(OSOF?&/B2SRW.EU&LJ^^
PZ?+G!M8EP]!!QB+5GS,%I)1ENI[9M,04)])R5*P>!%J?2(\0L[F<P-I6^<\,4S9]
PEG$@!@[[K3G2?-WUO433QR,>V)5#@HLGJ/47Y9 A]8F#Z 6RMLL?6:"TU2 WH<$V
P4^7Z;FB4@&-LCSKR]X=<55#)I3W3RK@+-"+G(:&"9E3<YJ 'USJPR;Y]4PIULI*.
P>DIJL]-+'C,&@:^$.?$=\O"8P H^'D'B%U-V.8FKRD,ONFVB]6QV\IO&X6E)LB?'
P\EWE>W6>*]0O@8I4"&'F4^XC6L!I'[<*,14!F-!69=G*+HC2/DAO,[%ME]-REC1?
P=5\DW<F99(AI=!6!4%?>B[M K-[,>[@[?J'NY&0/U6O;AQ]?OMI$ K#.1S_TG7/P
P<S'H,=W>;2_D4;31U2<OT6M$O(+#"1]Z50=F+P$$LA+,GV.,?VHT7_:%;3+(+Z1/
P6!4H]U[QB8."00VZ37@/"^,>X.>)!MQ?-UZ06:K"G5?,^#;M=Z-+F]JI^:IA;G[>
P]+>+/&:-MA]D^!U"= '>EDM.HP:_/VQNH]1,[(:P35+WG4&I&3[TPAC6*#K-5##M
PWIS>JY*.[H>$"6+DP,_LOL:#(+O8C]XUN#YO[UC,P=G(0#<O@" A72ADWT3"D2/D
P8!WS.0G/6!9[41)4?,#L%NJ"J->1[ _":[14/FWC,5E/H&),UYG):OS"C)""IE-B
PN)O9&UZZF[#9%';)MB8O(L_>B32TY,X.ZP!=UU<YD@M=YK*94,L!(EJT07(SHQN(
PVSXZ/#2^I+(1PU<G%.=VB]\3=0$06=+@.1?;T 84#[7IX0BB*#;6]_8$Z'[;6=U5
P=&9<0..3S@>!W,*MJR/&HOXJO["E?W(RE$2I0O@)'\V*UXD!1?BB_2-W91.;G=$9
PQ&@FE'"<X H1_&M%G,-$2-ZN_0';#,/F-L.OJL3:D+NP,"SO2=B3\!G>_%7:1J&G
P.6KNG'=B.U0R8"[/\(H48A7+9%VF/LNYTFK*7S=2!!\W7.*VJG:%VH2LY;I\6V_S
P]0;SX.7*Q+S<:U>PWZL.(3W(D_%2< =-DT$8'32G O7JBBICI*B"8>URIX4%9WPD
PSJUJ_.3;#M &@S+>'C,<JA]#ALOS&!H&I>%$P- X!1?!71 UP<XA_Z%)*UG*UUKX
PA<3EH,=<QOAO'$:61'4U[5EYC+HJEI07S!5T;\NXAN M:DNN/"0]#EB\VV3!8E;"
PZ0Y$K#(#M_M'=!@*;Q$':C,+M_H%6O.C"2 !8K=4Y&L8]'.EUT.8X-7(.[10(-:(
P+-_0U7F86\+5T)0^(WH$PQ!']GZ6L@RF2'AK8>E9@!'@CWN1'.]T3N+3%*,*AG"7
P_/!,[W?':N:)::IK4270(A1]I3.FR?&#3(>C[J!R(:@7WZ"BM .AYZ,SWG"?EP>P
P"/%.FCY,A3ITBBO9#:$P"P]S[M/9Z8"/.OG1/_!L)AT&*AF-Y,[A($%W)L_Z#%2(
P6\R6AS@6A>+7ECDH7+&9"G2\P@BL!P&7%I.^Z XD3LFFVDN9D$OB;<8!YAN5%TL6
P^L/U?X4@S7%6MM-KKIDY6SHB7+2A&^JT?V]*K.DD3QK/"K@Q3F\HIXB@9A_]V3A:
P:Q/'9HAE/EA7M=4=$,K@E3>SKU/.W D68\$XF;HI1SSTR:P>9:_N2EH;5[53"%9=
P\\<4/"5V%,- \U,.'&\&GQ3,N;4:<.L"7?X 4#N&Y &73/F.^A=KL6:WD*483G,6
P+,@A1+AB<NG06-2[:J$MU,K"5*664HL[CQ(]P>%4"+_.'>X'ZQW<<*(!H*'WSPIP
P:A(B,O$--P;: 1K[-F^"2X7AAP-1T-40C/RR2\\C"^X=B+&92AJP(C,JZ[B%QG2M
P^.NO R)^AS<:,(ETOFF:!V0(QPU?%XDD<@C%<;2!R@XA<@ZD5(6$QG3J=9@15.SC
P%=Y9+:@J72."-CZ$*AWWF($@-11Y#T\EK:4&<D7AG%\<9HKPC-$CFC&^>@[>"*[0
P5\]M/)4T.T0^6\69D?D3RH,H<.R_>(WB"O.J^>^:U@S,)&41L:"@4^^^)B-"F,1P
P!"?@@9<@BET@W"*2!?#6&*;>'8@ TIZ[_2\ZNJF(A#0J6/;9K.<-CD3W!T;,5<]>
PO^-VMB@&[&J.V)Y(B>A#V1O2@[L\ _4E83!J69^$V6>#0"##!'3ZB-*H9DQS\Q6Z
PFG#4X?',!6>F=C9DFOJ]20[R-"&#C<8F20!H-(LC^4RIPA/\_O,Q/@R^Y)* H 05
P%U5&)^?O7\R!W$W^G'^I =A+(*DPU!88I=]"H8@H%4/K"]]9*"DBD3-PD+/N 9.7
P .GA\.N:0UAQ92"L]I42MFA0)%_>SSX?+CKHJ!5'/,>U3%J-"Y;3-.N*U;-KXZLN
PY!RC;^J9IBYYP+!E[MVN+G:Y$\SR5 BAMEHN2!#YFA,=Z6+&81W%YX7@>/O0,K"@
P^$96/3 8'SD5^ZI#U=:GXL;E"3-_@55$EE/RN*(@E$)FXZZ Z2!@T"ZO"+^- =07
PDV6(39WPIK&13<J:Y"2X\S6N>\6YT@P3-YY"WSAWU;C%QN6(94B?H.)4?TXY^9V;
P7B.SZ-(S#]&.[,@'?>$_922B]7A,DFV4;J?10I:H3SCM1!C_D!U)6V;)[NL239ZF
P4[!%Y+&7\P!VS%ZR2QXAZ0QR%3/] [9[()";08$6FGD_:0P"UJ2B*1:;Z7GXAWUM
PW8E;LL,V_NR!@<#:<] 9(CX(:A2Q("#+EARXA>;D6&=M7Y06]L]8/3W=75VD8B&$
P"LW*(?<20&^8473I>!L7 "Z/C!T1&[+G>AQGJF>@P:]8%!GPDU@/*%\FK.?37II!
P1V4] EX49U'\6%W#D.(N%B4EB'O#[VK,*#9)F\W[2+!%KC>WLE)1NK7R<4B6!XEK
POKWR!]E4_1\>PJ;L"]D")]!K![3T25S/=']D\(S<QI>2T7-_ZZV#0OCYF7GVMB6+
PRH]P</?BD5>\B[-IUJX+>*,>;NV#W1[?U*(J!OZ$R$  WRM$FU/.RK) =HU#_1Z<
PQ<V2%@'9',GE?>B S< KK(;P '\&J:F]>)KIXA],#-KFON,?:450?G6;$FYA6/>)
PLRR!HE)C!,<H:O0@;?K(^F"O9<F!H),^ QU)HTV9A9OKU'Q>&#BD_T;8=@]*GI5:
PZGX;1+A>:9X&3YODU)J+><6-H3@*6-2?A "1K6%D-\$L;/\2-L[0&NGX2'RZ?YQ/
PJKFA/7 IBT_J/I=FOO4&*D1'*O(PW?41J@:9:,U^PU".#QFHX>LM>QS3U;*/7,3\
P:XHQ\(X4&%="$B-9K6W@NP9C!_=/-)&<NB6#ER ZN8^*&?KLT7^$VQW)PJI^-8^'
P&^_VE5OX,8_%X45]0MCH=:"*IH,0' KY1GN4UGV:+5W0!]TSO+8(M A6@[Y4F9,-
P^S.?UNM$$CZA7V7B_ [/6J<0;6%9[CFE6M!W'\O7Z^2VV)@6KJP,]$!S2]MT<8'9
`endprotected128

