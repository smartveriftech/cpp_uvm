// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
PIED--'S77*1!@?UV>HGDL"^E# BDCI0@/_N$U/U90X]H4<5VB#1/>[_3R!>L\7H(
P\4VTD#@+PREN_D]3<JOT.-*9<TQ)7I1)K$33AIN!KT=K7VT5A7ACV+B/OH,&<S=C
P(2 <X+>"<(M6:DCW$K]2WX7 #>_1KSM%[@0RT=]2QJ<FG?8KZ5_>FE!9P9B?OET$
P9OZ0&15 L5%(^GY)_R&R-I9^0MD<B8O@\L80&'%0HP[#CQOEE$UDMBF%R>K2CB)_
P#B'WSA5#W^O=P[1X;"7&/P&?$K\0&7KASMD$._0!DK<[E^:LURA7BJL8S@<K\IYE
`endprotected128

