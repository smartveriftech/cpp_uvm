// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`protected128
PL:QZF=!JSF&3TPH#08)3H_[,#EOJ ^1<G[##R2I9'_LY=\N+/3$44H$DS__U2[,V
P[H<%(&RC9'_)IL+9M.[T[D2HVRH5R[3);"+:#_/"BB4B,U/ S'AEB3 )[?6[_]H_
P"U$Q3E?*9JM DRR^"*C1"B\TKLY#=U.IU:,?,T"IV]C@XH76Y;>52)&/64%HI5M'
PLV&*/Z\HL%I*/:0SL'<-07^/S<-:5>?VBH$L+P.Q24DU,?[> G[>_ DU?FK*9)E=
PI'MF96Y1[\@FO',7WT#_K5ZOOIWH$%T3&_3HY<(VIQR%\ =\!\<$O_(V!J (1#M3
PY_U%OXW!)K9*1SY?:D6 "7KOQNC8S(! 3MI7! K*\SU7]#(8O1A":S,)BYF.+=UH
PK*-> .^L5\!YRZTL86!HB=''*"HI7G7NM>SOY&<+5AFV*WY60]ONMP,XG<FB8#AU
P G._./[[$NI]I>]>0:LGE"-*H 50M]P!03"9/-W*KCDX(D:8Q,0]ZKZ$-C\?Q:_"
P:BB)C0VZD#:*%$W!A6-PGS\F3@?P,/BW4W#G/H454UW%EW<JH.%$7]"LC?PD.1WL
P5AJ)V[) G_0UXLP?1<0EQF%_\[N'+:%O"@+;(XPGO"KK,/)].8CVC5,*G8QX"Y2M
P5QGMA#?ZB5F_?Y,8 P*3>P*"$8W6C1_\_]<M5BS(Q5:TN^ZBA_#^/6R= >XI!98+
P4KKW( L,I&:-I<II0TUD$8 $".7*W"/*>#J_VZ$C?WA8O\T[^6/RCX-@2GC?(<C%
P(.+_*_8RVLH8H+Y0E)&KY(N_;.52_#*+!K!';+1BK./2,PL:;#N+N66"*>7E6;@X
P0UQF2^!T-L\XG?#MIR1&RYES\_(="F%OOD)5N5BP&RQ=Q\"ECS*_%7B"NH8<3HXR
P.6//1;XKU?%>08!R:7$:2=3(>KP(B$7OS>$K5==$;7RR2T24S;FEQ6$)4SL,J:Z;
PC)$JN? #6:&W\]BEC_"-8K5U5:FW&>CJ^G N4JCK(NL]4IB6C;=]Z3<#6@<:D&A:
P<:BU1?$' H S>4C"+K8]&^B)9SSA@81==MT0'J7+=I&R^@X.\CZ!O5W_CC.9N9_M
PXPK'P)>,N$#)"PK#5&F@OM\,NH.<911'ORZ6%=K-!N,%/^QXE$#(KZ0.')55A[[0
PD!FY;906Z/GHJ#B>= JHKAXUE[FX_.H/HJ[Y!_ ._ZS&2Z4R>C<O="L&M'O]&S4N
PT-RV["/5&2OMU/OS%H.OKLSV+M]9,L6I>:+>.]:8^/U9313QN=TRQ$4]-)AH=D"<
PC<BEBM?R*)% 5_X)Y:AMG%MWMG)2C=FLE1!(.3NYGV)WSM"TOAU-;JHTND*JW& P
PR2Z%9N:R2N#PGBPVQ\.NRH#3PQ&EC)&2J$.6![+'D&&1O!?<XF:=;NRC>M,9;D1:
P3")6=PDX1L%5"&]! 6 YH)-E#PB&KZ5,^KXW)W-_GZ;\A'97BK ZF92D! +4RWEW
P\\N$<K&MU J#,0:]' 2""]9CF:\-*Z#+SCX>SCPDO<^9;7>6JE]8T.7;8>!6I/F9
PQPH&AU'URXB:X5[X]_V@!:ZPC%-$V1+I>]0]/FQLN'):7V@];]'*1_2KAX959O[N
P-Y+16-UPTFV66BF&(R42RP&1#,UT]&5]]JSBMS1MV789*1RYR*Z%53ZSQ"  MZ4Y
PR$LM3XEFE_7A'5&9HTD+F8%#S,2R[SF49MY)O$17J^QFWGQN>K=QH0X'(_2W@NBY
P/2:/E$DB_HJ%M/89&6.9MTT6H1=';"A3+^O\BG[]X*&E\0/2$;5-K7+W84EB&CNB
PR2-'-?$+<'\ X+1E.9+$XW*RL#*]72?EMD\5(8!0(LK3?SUA!-%)&U&.)E17,@+/
P2J-05%-Q.-T)G@6J,WY9_9/TU>&/75WK$SKUAT'?I%I.=,$A(=L<M?U9:DR&PA9=
P^O#WKBJ>.Q222Z8RDZ(..ICN2F>?&8>DT._MS*W (*X^/0<#WID+,EU6E'3^+'; 
P^[4I.Y*H^0DQT@=C2GNJ>0SOH$P2;@4CWFTU6<C,DOFQIV7.')4J-)69OX1$C0I.
PF$+8$Q:'N*4E?,L9/1G"2#;^LU9X]^S<^0^+OZ'<7XBFA4+;UI&DI2B#V.[:T>WZ
PJ)U\X?QX;=9GS?RY0#MOJ*>Y?D_D5OZT%:CY4KY'S#38C5CA'JNMO*#8WC.$6>I9
P(RK4?$R6PH'%QR=:.PIK-[\T??/ROK-EH\%[B8$HHW#;41*5:60Z_>47>5]R LGC
P"R41J?VC,3L&^&X8;]U_B".04Z5<SJ#05\B?Z:O[UOCXV+4Y-OBAF2T5523UAY79
PE)>T#N&PW2F966B *YVQCT&$+7B'+[@35MO7W:Z=1&//P+F; .N>9GL7OSS7TD'Q
PK77K. &*'4BF7[*T>H#VW: 40/TK&O%T\S_S$^-+M[A.4C\MZ<AG8"7L(G5\V8-]
PU\^ #0;0HEBM5N<I8XH0P<R'+>$<L3$D>5PA]0HR9I5L>C3C;L[T&^F8'O)T;48[
P@BX,7]"UQ4O=B^N24++-N)B8[1Z_M:..8$V0JL;B G&J41_;*6OO<+>\MZ[\T"Z#
POPQ":-F?8P#EJ;C4[RRS7F<4'V=9%94_R+/>2AOQ6XZSW<DP3:WPC#I!?-L*N'<!
P*GZ:E6>*&2U!;RN<^\**@K%0XRP$?C MQ6WEKG"$\I^HE$+&\)4( SAZ36:1>F,7
PQN(SU][QG[AL1__1KQ2F$4DR5J8E,C'*"?,P%Q:'ROW_[0BXW4(CSI'*<-A)"=()
PV#!#=FK60F+3U*B8@EA![P+/Z'$5^%X3W2%.Z/*96F56WG/3^KQ(FBXH^K[<T.NG
P."W]R,8 86HT:P! Y:GP.3[!SHBDP/X%$!P;K3.- _U)_3:91OZMAF7>F5&^+0>0
P=Q8R"4-G0BW="H)2/24#1>U@IC^[=7BT5@ ,,NK VG&MQ8IN59@<"#ZT#R^"Q<HC
PD,Q<>1H%P^U0)#W(D^()XAIW(*XR0F(4O<<A3_@4P_.)30*KB:GW6X>GTWXV'P"#
P4@\DAJLWT2&;FKN#O#+K]]E11K&PX)$4-ZN/:$WLF0'YO]Q G[&S\PR^EP@.3I O
P-Y.Y?,G\4U#W[Q\2W*:\=^/?PAVG$F<ZI73*RZ5QH"Z]7"2KJ<=/\^C-+[.VHTR.
P-?8:#M]52BAM!70]=0,L %GB)(0:N,%]-T6>?93XL.?N'CA>::BFTG'R=TB;[MS:
P\A_=*$Z_H6= YY2>42NV":ID(D8PE_Y-9[L1DGTWLK\;)&%T;W2&$K=X"M 4U@9[
PH#CY31MH$F=GM1ZS6E$^SL;>]T7QXD79:9NAU!<:4);T?&;HM_^5&;F>I=^/%/'G
PUJ_35(SBU1?>T%,<SXG'?+K[S*-H>0ZR!H<]K.D-YVO@VHOE6:[603G[*\3\:4T_
PLA),,NFS([DVAQ3D*%9)!%+$6F "Y:4!,;G8O&"C,^/[=<]9PD@G$'K]S#@W]_@@
P9LY[@:P5=]:E0[=+S^4:&8OLU;O2XVA?_<WH\[#63VHX* KJ<QI9ABL6.QJ6I=F#
P?IX*<W UD8@UE6'3U'!VIYEC;NSH?_2N?&W_BWX.C9%W9,YH.D[)MCK(.GWSK#%2
PEO_%N,K3^>K<'%@H\U14NH0@364DZ6S\Q5I1#W[9->MQN^'SEJK/?R)AUS^_WYQ$
PB6K>KC!.'B?;J\_!:A0'0A[[EPG_I/_![YMP;P.G+*D0K^MM]+K"Y.4\9+S/45-T
PN;I$MO4_5+I\PV=U4*4^?/:]=G.J %Y7/,7KVO XB!=S6;EC438>$8.WCJ=F$3*L
PEU#80P^2CZ'(^YPDY)D:<A"]P:KD:ELK(H)'.2F"4^[>6 SK='.Y_$T:"KY1O+-.
P ,>0W.',.IZ#S^R)!WL)$LQV=F;DC<:SB+A."81;L\7SS9PH<4NA"06/Z-.(>9@'
P)7'NCI\I='X]#0=,5LS*F'@UMN0@ .QP!/\OSROIMVA5(XBV3F1T,5O$#^Y&%"DY
P%*8C+\K29FL*< %X*@#8J$7]CRYS3#_6F()--+WXGR0"^XF)_EEX(P^T^)R5I'C.
P=U)X)7MV6G(&;VAM!_:Y>$"S;Q>@LY@X99&G3NN3(\3=Q%EGDU;GF2RGTA[LW=/;
P/38BK/(,)%+7[J'LKA\NL9;_+H?>^CYCG*+&^H#Y'1*7#<PF,*0GWMC9H"F=#*GZ
PG20"]=&?$M^8DBBW)-6?;[H@(/%RSLY+C3Y@17SC"/D*/#M8&0U,9-9\ @U,*0R$
P!  J<%1$AS,  ^$QQ&S=A,[;[FB5T;I"+=VTJH]O3245?W4.&/'CM69C9X!PK*'B
P@'4>$"H=AP7T)X$8R]/HI##;0%_ME3Z9VG?3O2\77L?9<&",3X*;_/O/MS5F:?^@
PV& 7ZJ.<W E5_591&N8)C&H4+KX_]Z3@K*O%JD&@6J?A^&Y^TM8]04"5CU)C(:;]
PE K9)><U7&+O'/.N;0+KH3X+:VC32%:AW\&Y$PB%1-N9\[9#G*V!FP#AJ:R*W&ID
P=><4$V;BUK^J$#4#:.:^(KZN.N\\XA\^CF(C2S3[F^FZR>R;J_,$'@K^'T@GB)K7
P<%7&]FVG:C4/ WW"2E0G1F+W (QC><T] B7EEX641<<_R<; T[23&^9^[>7GE@0R
PNO/L+F5S8;XLF4!LD=LM8#/>)SMKGEUQ+/#C9WU6UD54K*$".\5Q<E*,?'2._NVB
P6O)-7)@U+;HU,#@Z>EUNJV+$K!A_#>?/T\-,8<N6=QW:"'RSV)\M4EW= (C45)4>
P%LP(9:%WFW@QL'R=9[..8EVJF_^(/YF!-YK$BC89FC(J_[7FSJS(E^\ _[5<JL&<
P0X^T)<V7KOH1MIU[#HI$*.A&BR1&&U_D :_@<-)I"VP*6W/7\EJN)DO8%9[KY=T[
P95\XBS+1[>V!J&O^6QF]9'%F*/9-)FM0T"]A>ZF[JD]*=LC>_0X([J>9HV5J\4#L
PCB?[CSR5TN2@#Q,#^]W/%Z>SNY)3KK5;GE3LQ@QED$]<>ROI=+X4J<7X9RQ0CWN0
P="0LK&;Y#(]G8<HK4IN[X(Y.Z'KMF(8QBXKT^4O#HIK20^YD)G1\Z8]-".V>]"#7
P81Y\JZ/=I_$3P)VS&"^FE; '1BH]& <O>;?]SA7KZZX55UWY4 NO,F ^RLD+ATS9
P,%9&9]"XIH/.NX?E=/5.F-><"+,5?$_K$@(M9D?^B=QB13H_*%4TF5Y#_A3R#*DF
PZ/NUP P!.^=E9+*IER$=WX(M#%$%XCF4F&AW#E. *<3@$;I@,KK,XO7D_5<*F%WP
PI3M,<[RCBPE>2@@.5X&Q 7L $QB8>QAW4*N<03=$Z?L/H$0+-$VD.$AI=]'C_K*+
PUHP/U]0G&HZ/517X_++<9B@T=GK8<Q*)O&+K-?S=];D!]'FC^ BT;8_7BF;.UC1L
P19_>9Y+)4A"[JFD\3['Z[SU"!Y*\-=Q5"I=1/,])=J TMHJ82DJIBZ@QY'T[E/U4
PX+.Q2"M)U.4P3J]/-7>^:T$4H4SJDK\$Y<=7E7QX>UMW[Z8L?2D:]^V*PY.E3#>X
PG5O5!L'!P-0M9YI0<FU$%J/XREJ&]GGXB[=N9T?P0RHQ4IMED3V<:E*DR0U%!/>Q
P&P(DK^3V1&(N>)W!TR;XL4_",<3ELFH%TEGN:<D< L4?LV/ $X5KQJ1"O9;VCJ3\
P7ZVBCQ+,GYN!U^.K^U(I"L\*MKSU_,+_1&3LH>BB6@RB>&3Q"?1>T+Y84P<Y)$9<
P,MH6&ML_= N7Q!7"+ABGQ+P0+WRS$DN@4[QDE@+_*,]?#4Q1-YR"]]=$HPM81W-^
PK#9T#]6IO,NDOTIFBEIQN:_40X.(B"NF'[Y.7_L@S8AXU@@%XI? DL56:ETQ$8M3
P='F1VP#QV[R;-SRT[@CX(:N32F6,NWFV5:'9&5TKTU%XLIN+5))>FI?*H0W^^7S,
P%/C_NBWW!:06U:3-A_;)YC)TYHF14(L:.2[NJ"V*4M)T/;"Q\6.^-'0PC?_I>[@R
PO1*;Y+@V.P<TDCACOY5M'B<+&PD1$SD%%OT>>COC[EJ/D6$Y:VQ'?N C6B4=RS*$
P;#>;]R^(29@!/7PEG/K(58F"Q4G+62FD[<7@'Q%M"0IHT1ZSH/Y*.7>GOAGV!5R"
POCP.HYG3\Z^Q1'@Y-NU7Q)D"K6JF !1*9<H+/O1RT5'?G#LZPYG!F)8\X!#3-?E!
PMC;A0^C7X!8[6T /[9!?)37R>!S@U#C>@ _?,*;5@SVUG\0SGG&J.(5E]5!]8&D\
PD)-O[K[)N(QA8QV(+,+\FQO SD0DY>=O_V5#H[;[3O0/;B3JK&+P)/\&XV\3[-HM
P8//MW(M5(4$@9X-"1+ZF_U:-<L/#E1SDO$3NM &1(%/ES#;3_O,1R]1"GE9AC'^T
PDMEV"G#]+XFC(8>C8HCA'G,A6'#_Z@"<**IZNY-5AUW2K8&I2\O;1:F(SD2N\1CT
PZ>8ZCK:R5!WH_A(LQOM(&:Q%=9TM"D)C0"[.)S@;0<]TR_.S6HADMY9D^:ALTK><
P;"^A(:2O]ZJDA5KS"_G."!F4"R5Y13[KN1BH8MQ;+PF)6_/$-"NZF&T)$)AG=%9K
PU%06&S#P^C!=#!8S_,:GP7+XO8GVM^Q#1O&$''JPYV;KLP55$BV0^O!%96M_FJ8@
P2!&O J\QJPYOXASVJA*(%"9D$.OH5&X/#MS@H/7<B!A7_C]/B2\B&AS>ZI:>,QP_
P/FC"+V+D#EF_B ,*K$M,GR0_-\)[7!(OD)ZLNL%)B=U.(QK"VZZ6/()$9>-NI^:1
P<FGK*+@R$2PX%$^YA<!Z3,(';*04T@5'_2S'[>%M\_;!E2?+_R*$E=UQ>?:LK[<>
P0235( G(G\A1@2$N!XJ!&H[,&A .\6:Z6ZW/2E.582D#L5GC![NU/*=@K9&]BZ,S
PHQKZM9@?89_+C?4N#;'A9MK#OC;S-;XK1>I3[, 9].UM(]L!O[C02#(<P@DO9XF^
P"F^R_*Z$U4@)K!S[%EDJM,<3(1JQ1=FE*#%.>R(V&KX<P8/-E#YX!#[FLMN['BQ:
P89]6=8:Y2M2S?4J^W9"1:('OW,1=_N>%YJL)]Y=2#AY%F&8VR(O0=K?#6,D=\Q28
P 1E+5HK4-:2-*^"D5D=7 H?R]NDM*1PT,)5V\RCL%Q=R<^XV[4"WZO&#+Z-!"^9;
PT<B+M8$9J$&X]X20^'2TI!/ZF.!B)T(#=\L>ZP[)0[B/1MRJQ$T$=7BR5B@K]AE!
PZ.K4-L6G42PC6& \'17":C1/8MQ0?$-FLT+$A!'GB\B5"L+;)VFNU4L_NEHM:6?Q
PG>@$_\GGE;Z1A")A[CLS"V6A O=(P-P*:_\<.=^A(XW>1BQ<=O[B+@:>3>R^9RLD
P(;Y]=.*B#(??V69XQ"BE'RG_N?A@= XI +\ODAVF04)]KXE-+'0$3Y6.X8L#HW&*
P5S*&@#/7MDFO^ISY"8G;?.JW=EFS@)+6AFA,]34E-N':D*1[T&G ;J],\!1[,*NS
`endprotected128

