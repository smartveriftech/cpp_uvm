// Copyright (c) 2025-2035 Smart Verification Technology Corporation (智验科技)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// File: uvm_dpi_common_defines.svh

`protected128
PNXXYT 6UT[+5=2GX&".[\BIZ)E2&K[=(8VT]D+C3BBT>WUR":K>MN)XS+'6\'ENE
P5SCA0ZA@:RCGGJ#QGIXR%>/ITHO?"7G\I5*_ #NC[+4^<L,]HJEXV#L2<Q\U,$$.
P,K!?^55>Q'KE6T/-X%C9*9M[XL_'$J\1=S>NI1Z$62_ DP3^NXA(Q H1Z/N2KDO4
PM*I'*>GB< HD;$#O]H49BX!WA":9_*1E:7'CF;^>"_::B4MS&'YP<\/X1-EK!W<1
PN,JI$ H9F,+^R#GM"K5??Q]N*Q1(?EAK5GX[83IFSS-*3[Q)^W9IA4S0/%Q>8[TR
PAMS941\D)ZS:H?7WR61GC4M;3]-HNHXJ/6+0^%I?M/]V7Z)H-M9X\"SIQ:(AHH#4
P_")/]9)"5ME63@,:$*J@T%EWGOXCVSQ K<8FMTA0V=O5BEO(@+_.E4O37%0I'6.]
PZ_B>0T?;;;:27/4BD#N**YE);2I/+3@:7I;84@S=XR]MX[;P9'6),KU$(Q96@04U
PJ(J,G\KQ=N16OT@4>M0&O?]?!6I^T2$OZ[QC_8:? :-(178JWF6G$%W52F;V5:(S
PH9,%-.O*6"YF3R%HT18\+IK+3[&/-:2;^/@>.-\13#QU^<;U!Z;&/+*2$<TO!>CJ
P:.0J5&\?I0]4\<_TD;09JT;*DD:- 1/Y*(D:':$0/5/<OMYDEW(:?D#?C:U2VKHE
P,8:L6J&%/_!L76SB ;ITQ^+B"\Q1FH HZT[)\*AZ8.B&7:N\'9"VH%W1_[0%B0UO
PS*7&>5X:R=-ZM\@KX;4/%->$]L%5BC*#H]S9S&OW%.5\)HU8\QXEO9]VY_?U"3LQ
P3.*E^1I1C, S"ML54VYO;_C_!]F"W#+/+SC[IV0O/'R2:FP.>PH?VTXEAB5(?'DW
P&UZ7AUU, C[MK[$CWX4-\7QD=[>D:?VY/+-MU/"!2XD/N$0FNM>XB%FR(,X0RGDK
P@.R5O_V^I0#/&\J'5U!2*^[?:V9%)].8]N3=I-K!1D^F4@+3XFP_TY'"/3A8$+E>
PYV<)DV^A,5SS^<XO.'D>IPP8QF9?Y9W[0^-%5 4 56@V[7U6Y2-B6L=1 $T-3W\Z
P2H,FSE\5=[[3*MW7*K;<PTX-W5+"U=S?@?3/ZGA=H )X>^&'+\VM4>3]3W^:LX!M
P!+*O'&<NNIH8;6:H["E2DNQD&H3GG515.;^4W$//$=Y&EW5_E(ZT-':C%B>DYJRE
P:C<.,+HR#;R(2"XMLP'OXXUOPH87F.<XGCW4R9Q9\D%WD@Z[7PQ,4DOJ(Q4@\2_6
P0ZJV6;,%7UBU _7/-R*O0S83EU5E]^KJ8K!-[1[X?-0<\B2J7IB"* ]' &F?$H.9
PH"<*Y[VR@>P,O'+/DO#01X#K]+#S]1?!*]IIS]].)_?Z,4,%$Q<<K3T]"%'SFGWV
PY'\5_NH#PU"ZN,;@MRQ>U8K/,QS!&?/P:J (=SA-YJOIL!@=<4$'75D;#LM9?+P!
P5#>N6&3W<Y.UT7PL8#FE^UQ':6$:]&O YZ%)>_8GE0\"^4/CWS8]MJ4B_0KA+/?/
P)B#&-'UT/;GF&V8 :.[&7 OM"J2<U]2HKV&?KYV/6-S75_1//Z/-<-#PB>AFD5A 
P %F_CC(3"JK6NQ$K?GUJ&IR=:N2,-#AHY/#;YJ""L_G-^Y%XEH2>G-0+ $( _<$G
PN2FSK?QHX!9<D+-;.N.^B212NZ@=#1<EC=UM%%<ZD^IU"/8'_AZ QC_R2W;57OS(
P08P><+!JE$\85WZ98(W(TR.3Y^7A[)T80=@*HE3*:Z]6)UF':DJA8?I[.@C@Y23O
PUBH\<<11YY9@[<;3@^Q*IM5[<;W/'YB=AH;/9%:ME1 \XB/^JFZFCP=OJ&6^UQZL
P;/MV:QX;2S L*<LLDY%Q;UJ73 -*\8'>Z+$.&[VF8F9@2[?5^5ZP^O%LG9C[BY2)
P!Y"[\X+UX>]Q;:806T;L^+%$9Y%U-4]J+@.](/I*$[L7#XY7*1B[&#^$XLL)NE%*
PA-(GC?0M&WYF&X1C('BHM_IZ@#ZRUXRT/#>I]MA%_KL.N5T2[:.;TE)+YE"^?R;(
PN T?TBM?L7K21B,(E7#A7SLY7P/\^E_SF%#C1.KT5;"?1EO*C!!'>[R%B5=&>.[C
POGRND8-5_;C,#I"/]U-,>LX_9$J^#375=]H R ]BG$U:'"K13B#J5_CD"9]S&!H"
PO-@TU(S9S911Z)":!>%SM[BC.SP/P8F,L;;_)J_8;!=?#[+?#X2RPU'5^:#8:E?!
P7ZPL@8C+72"GOKS(PZKM5)RV+/*@I2 /\99BKB&\"9*::!<">U4:C^+%@:6B9%.V
PVAZ624;Q""(H86-L8>3$3C5Y<7M8;*E_87_MK%EQ+L,_/FY3']7W6)J.L8@$^)E^
P^W(3YRNPM$9J,Q_J"&A=*#G8S,: G&WBV )K=7T+U?%5^NY'^XY3*/W%A(Q2:UOA
P-R$";4@Y6>/Q$+?%:%O]O7.&X8P])+[>.!"*$UF(!##"7PPJZ2=1,*D6;&/%_/[F
P<5[)9LNS$;\BVUG1?M'KLD^$%41OK)I::V;)99+ <3,@*D$-/\?36#JOX\MD][JY
P /X/ ?DU:2S\/=2DDK#BLGPYW*?Y\RD)G,)>\TC[; _(_8AY=.1/LM]_UXE4W1>U
P8,NZA,T0QRD/%+I!(X A3WTV+[^TMR.[$@V;G^M=IYEC[^4-BB)\AFQ/L*@K%G6@
P ]T_H+CI,)C+CYCY>W.5\4I[9W?\S(YMP6E'GA/QMOK/*?MV*KHIKG _E/I0/&$<
P\V*,>]=S4;\,2QLDPAO&39(BJ?I$/2Q5'SF^K$J'^VGF;\MG/;=GS*P3-0^1=0U8
PIJ0GRXM"(2TL&W)Z "E1^@'I>MHQDQ\W)OE+2*=4$=##K%O U68RDH:%[40I6;GK
PC)!0AS#02H1:,J2?ZID[SOP@&)BHZ0.G\8MPT 5*!2K/VZU]^K@8XH .71\?FF_?
P8X,(C>SCZHY3?M=3*"*2'GQE9K0?0;IGD:4(,6(+GTR*4<A4_C6E5;#3+$([^4%@
PA: /0*2TPCS/AXI@_FLYMP)Q^G>\/3;YRL9; JP<4N<6Z5YJO#QX/R5Y-"35WB:X
PAV X@W;2E/T_4RUX;\3#I@?8JC6AE>HSHCEXZXH3M>U708NDG,07N64=W90FV!<X
PO ' 6=]B7N<.L&I33H6G1M?">)("%[XD+"R9-4I_.&]$"46RIZP$[$CFK!*R8M_.
P5AP&C7,::*7C("?'-F.G:V3K:+EE-X(TI!Z9MJ'@W=<M2#I!)9,<[_6!0\O8)8YL
P?1T*S]MW@J@9+VXEI937G.Z51K(8BB5I<T$TQ]&1.#73(%*5(?:9Z'YZ>FTL^N7V
PY$!D"@AH.==.@!BZ]9_<BBYU<66Y4EFW_$0?'VBHT-_T=!)FS\JYU))<E\OTO5*9
P.N@CH4!Y])!#LC,#KKY+#H/\BDL,\H>GK<_T*$V?3W*$.;7TW>'5@>2G"[1B$'CC
P_A0F?)M^'F=^+IGOKNN 1PLA^^Z7T )1QI=9_L+G(:M2,!&F8O=\Z0EROJY25U9T
P)%D-XI1/#@6,!8RMD(H+/]IJ,]782<3D8.L_Y.K&H!UQ]355!G+XK.&"X>\IX#:V
P^6H9.XF1FF_362SE/4+.D _%U(!JF$ =/M-[KW1#2D$WW[3-SS]@Q!@S74ZR(+OB
PZ4=#Q0,<H9_.9Y\4UV^S/CYH^LBJ(ZF.Z*U'?,)@HF-0S?K#UIWJ<PDJ!=ECF\H0
P8W-E7+-TA)C'L-J6 R\Q__IZ$4K0&73MJ1823ICY[CXVNT?=J)'&9/^\CCNNG4W2
P[)L^(HN;&B+\FI75$3ZK1;%[D]LD65>O+#=!:3>S !#I#AIH,ZD5Z<GKZ^?Z)J]S
PUE7Q#3KH$LXB5X(J9'M&#TLQY2#[-;]#5+G:]8+&O3WYGI4+K'F&#VBSE?NBD_[*
PTQY9^?4RU'&'U]@#:C-(,VZ6XU)I;W5G 2L^;;$(O<)I>Q'QZDDQR+)H.5J]"Z8<
PL#\=;P2?R/&^(X=?KQ\K5=CV<A\G$K&JOPX998'7"0+%QD%_>DN@*Q<SR_ &3=HG
P"=Q5"H8G_A144/.,>='+47!6[@YE"B;Q1T@,3<?GM2--\E8_M"ZA!!NULZN*Z6_S
P?\NTXO)^)6CZ5)0>:OUB>V5O[8^:B4HJ)1KU!%#_3@$-?0("G9+"/WJ[C6)ST8IJ
PE>.*&F.2(2AMZHP)QU!?HREO*I8HU]YNLYV]8G)X$EI^JGEHU+4K2767;9T%R5=J
`endprotected128

